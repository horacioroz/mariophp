            �     (       @         �                 �    �  ��    � � �  �� ��� ��� �    �   �    � � �  �� ��� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� �@� �@� �@� �@� @@�  @� � � � � � � � � @ �   � ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� �@� �@� �@� �@� @@�  @� � � � � � � � � @ �   � ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� �@� �@� �@� �@� @@�  @� � � � � � � � � @ �   � ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� �@� �@� �@� �@� @@�  @� � � � � � � � � @ �   � ��@ ��@ ��@ ��@ @�@  �@ ��@ ��@ ��@ ��@ @�@  �@ ��@ ��@ ��@ ��@ @�@  �@ ��@ ��@ ��@ ��@ @�@  �@ �@@ �@@ �@@ �@@ @@@  @@ � @ � @ � @ � @ @ @   @ ��  ��  ��  ��  @�   �  ��  ��  ��  ��  @�   �  ��  ��  ��  ��  @�   �  ��  ��  ��  ��  @�   �  �@  �@  �@  �@  @@   @  �   �   �   �   @                                                                                                                                                    	 				 		                               		 		                                        

 

                   hhh            hhh                     		 	             								        								   hhh				 hhh								                                                                                                                                                                      Cadlink Version 1.0
 �P�B���*N�P1�iP�)�9\�l#fS�y�D7n�lN�f=�r���p�lj[,@�LLk,�2�ِ1���z ������(�!fNZ��u�KV�Y���I�>����&&A|5j��'A��IT� q��I�WK��E¢�j��&.��v8fȘ�M����C�A���$C����z�Yϸ��@p�q�(�&ޫ疓h_Ak��fըُ�'֠	�&i�hL\�{�
0����������Nv7���h��j�$�78�V-�h���Ĥ���nb�7~�I�~��?�T��wiN�8�#h@�҅�Ԁ#B1�Y��A�(X�y�HC&R��'F3�$��}�ƒ9�b���3�(ps��$1��L�$	mk�x���+���&����#��KK̙�ӌh���ZP�$�gJ�d��������H�q�=��&>�&c
")���$+ƓHR��c]�c�7j�c���I�ȑc��d8��_M4+�D�[�Jq\��O�����I�+4pb��W�W	�W�"i�`��H��#��$��K���IQ��d*#(R�XY;.h��aæn6��ѡ&.�����Ŷ0�Y2fĘY�Z�(5���F����.�X^���z��U���K�.^���Q�\��9Q�e!��rUs��,�[����r�W~�oh�<�.!A����X�pS��v�T��T��ӄI��[��'S�V�zj��Q�4���.�ZV���Z0�뫩�B0�0U�����tђ��K���%3r��6���lba<Z�ɬ��%�.����87-r	9���))FLN�f��]+3���X�%�w҂A�N���ں!�Q8�r�.���K��RF��J��钳i�ͨ1�3d�d5�,��Z���mJ��;]WEM��W�w6r֬Sm�<��Ͱ&�F�
_�fSr؀!sf,�4�%l�0r��iu��R�Yrd�Tk�.l�<� �%�a���z-8���p����6�P&��]�F΁s+0��W�âps�Q7��Ⱥ+��U63%�M�As��qS��N�Qcf���.Y��v�_hɸt�.����\O9b��"ݦ����疜�v�ג%.f�/<�1]�把�1KXLua��dU�5[�Nd�5뱬Y���a+�%��b�/6]2�z&mv�©%��ΒY�ݨ���m��:k�T�9�扫Yh�����Ÿ��R�~K�̝�`��n��5}��\��K2���r�*�����-?�M��f�dfu��uY�q.�������v�{�)Y��}f.�M�-��;��w3͙,��$f#S��n������":U/<5�{g�TX��f��.�̲_�S��j�,,j�p9e�5�M-a2p���.Q3
���.�|���͙v��.��A�3�q��SW�g�����՜�]qү4h���c��a3ݦK�9\¹M�USm��W�-�ih�d���A�v� ��.Y�W�u��~�����bu	���3m�dڦݓ`%6��f�)���,v7]��XLȊ�I(�����4���iI��	i�sv��Ŭ�%XRU���̰M�V��?�^r��J���uIz��.9V��ű��U-Y��q�u�ڞ�nb����8�WdќdŬ)���؅�d�`��IQx_gS��(��ب	K�0F+Y�'���m�M8�F(l[�*+L�!��-m* 4r������{�^/N��qe�_r����2�R�B��f�M��f�<�J�!1���[rO�܎�)���YX�;g&ƅp֒���̗�PqJ��dҕ@�h37��R��%kg����SK����J1p�σ��I�F�
+F7%f��x.k��q��嵒S�:�6�Vb�9ٻd�fS�u^�
2bȜ��$�,L+�����1���Z��9�W������\KM�Ĺ�������hƱA��hԼ�"�T�3�3�bh����x��R�@�s/䬀Zr��p�Y�d=��j��t	��n���狜p�S�P#�#����8�T�K�'��M�I�rY���/6��$1��Ui�l�x;ŘIps���S��k�E�}x�
���@��԰/]x���ͦ�?���;G���rXtsb�AShw�5b*�]@p��f��H	[a)Y���r�����`3ǐ�����S��FM�B#�,�+��+��䱸�M�����\v7�o�%�VX��X\oXljɒ��AN)!#��ߺ3��l}�y���T��\�p�/7�_X��0}�^��Bb�Wa-9�����bզS��:͐�ʌ(�v6���f����k��Z�8h�-'-�]v1���L�
�D͡e�ۘ(93N{7�)��\�ZTfR��: �*9���,�k���j����m~%�~��i��0I�(���K�\��!��"K���b+��E�Xdj��sX:��6����F֤9�b�X�koF�B�S���#f੖l̩8�&��qBj;P�PAJ�T�E��r-KH���Td& 9n"V�᲌�:,/Z�4��%lN��-��LX҆�0Z�b沙��搿^llcaۺ����`�13hЄ%m��\�e�Ȏ?5p6���eU�vո9ع	O��TE�ayx���^Ɛ� �����4��23��Z6nؠ����+�~�6��A@�r^���3k��M��:7̯��%�n�t�+W0d�L'����p��iI�VXKȰYa�x�AM۳T�,եhf3y�y�O0h�M�-�L�!��17py�Y�Gn������czҍ�v�b�'�Vf�Č2h���]�lF2���d��;�pU\mb�_d7l�O��\хfy�ck�%����j+L�ԍ0v���H���u�%f��CK�g�F���1j"6]����·8�զ�y�Y��p��Ԓ�q�[W9gpҍ�vɢ�r�Y��j�2ؼ��u��T7�GΉ��E��d����9zrv�`{��yA�ia�A�@l���q!\u]�Pn�ȁ�
1l�e[�9��<y�.��1��2DS�h���U��p�䐾�����57g3����᫫��Ir-#���f٪9��t���1�'T�f���%��+�<����fg��Bnɜ���S�LUa,�%W�_b:�X��z��T}����\�������.U
5�y1+}a6���[��M�Ir=|u��ƞ���a�L� +8U�QL�,S9ۭ�����S8�m,�`s��_���8-���mr�b�[a)9
6&瘁��/�e��!��^��R>�ߊ�f͔�����U+d%�ib���.���j.�������@��j��.����e��o�.ލ-�"�U8��T��D��f�~8�1f�6+���/5��0�̚�P>\��d�����M�l�͵\C0l*���3κ�l�b��Y�˰�p�H�XG6�uD3�|�±Ln�A{�c #\��7�\6�t�9^�y��¢:�^B�������6l�d�Ĝ�`]������|���t>���MEa,�2���A��n���6��5]����s�j�%���jN<4d��"l�Q6�0����mZ��g�X�%���7���f���Tu���P4�H�XJ��๹�J�E���/լ��D�Ip&��]"�ޯ8+L���]����3\�\˥gە�SY�F�1hY�����h~�k=ɐن�w,\+8u#��]Bf�l)������7��Fƍ���%�x�(�iEVl�)�b�N�3�qn|�fm��n�����K��
_Q1�m��@u���l�2U	4g��76lr�%d��k��M-Y`ݬ��Vl���8jV�b>�w�$���.��K~�
ߦdm.�!�����Y���}6pVINWܢE}����R��k"��-�6�ͳ���>��&I���0��Y�E-g����%��"!s0�O��Z��-������vm7�f�co�!�6\�KNl7���|o0,i��d��y��&fc�V�rp&mʆ�v�f��ã���)`���}ֹ�%p�����9_�y�'s�9��d��*�4��j�a�|ɰ��9�n���%h���dԈ#�<&C����9���M�l��?D�Y9lj�R��f�\m6nj����G[�j��q��b��.A���d��1E0�*7C`4]��ߦMoPL-y,7���������,�l.���3���Z�E�t#l�]��΍×���Ri�\8�6�L��a���5f�����;��d���	g,f�<:�N5"-T�rsC&�F�
�Dβ�
�x�5���-1`�T{��!c��s��XZ0ϩ��Ͷl�T��ҭ�m*.����Kg�U�
5���]�Ĭ�;�`�>�M����sy�Ԓe�*d���i�݌�H�l�L-9�E�a��a�/\K_L�y��j��_��Q5���<Ts@8�����e��!sJ��{ ʌ�h�oJ�M��mxa�[�M���:L���l[�f�;�t������=�|����w�d}���~��)6�$����)94-��EN��*��x�����K��gÆM��uDs���9��i�/�`Na8hZ�{#7}M�M�v=�0+`9Ġ \����O�u�SYt�ro�Ս���9B̈96��2߂s�
�%�6V�k�t6C��(&����u�ao1��x���s�ج��k��t���p~��X����j"3d���{���3�R7�u1���.Y�ͻ�Q[�qS�/<G��_�����#�dS�9�6�f�h�/1�`�Y~k�Dn&^M5td�>9	�ca�,��5�<7]�LԀy����.Y-4g�2�M-AÆ̹��^�\X����L1o��2����$N��[�%j.�i"g��4����>��Yɴa+�%m2���|�lN2r�Z\1I%�VXJΥ_G��)5��A�	1���-�?�f*��pNZ8끦�p��W�%ip_�f���cc���7m�W����oZ���4�ϻS����m�KĬ��3fK3p�n~�nY����T+{����PL->a�Ҹ�%�� t��N�n����\1S��t�7��s��L��������A�%hZ��2j�Ёi�`�{=7�fMc8��Zp�]_2g0nj���}m����^*�;/��2n����T����K��9K	0+��zl2	�a+�%��dɬ@4����}��)]r��/��B4�.⸩%�˦�Y�CS�S���~�SC&A�0֒��ߌ�`9˩R�9`��-���M-yv7�p�w���,������
7�U3�;�p�f����ĸ��Zr8��p�Tʿz�EvE�钍lx��Y��aS�u��!�28Ս���w���D`s�.�ͰI���Zr*�+��u�l�$g��M���Y��\|h�C#�1k{f����%������,o5�p�ȰI@Nk�r��^�_Z�5��C���IK�_H`V�LS���c��Y�RrB.n0Ǌ�
j�n��2bb8��R� �9��jj�a�z>��S-S1�8�+�ݤ+�*l��&7�x�.�F�ϫ�8C��L��*,%f����`���``���z�eaOV9r�g���ɬ�������`�T=��O%g]�1.������=fV����%��(:U�db��ٲH�\0�S29�;�S�9tl��[T-D7�nE�,�_Pc�Wa�T1b���l�u��۽䖃2h
�on�wլ7��ɼ0߰uX���41d��i�.�d��Z/��Ǚ�֒{�f�o�.�"���rd��)�/�Љl����Z��J��I�A�ȓ#�&R���7���a+�%+�ᘘ�������5$S%z����k��J����$�ۘf��
:����BFN�J��X���Ip&�����q��Yb�j��̾���̹2f���(�c)��s�W7���u��k�M����
=M�$P��Z����W�T,0�f��T{���f]���T�ɹU�ʩ%�|�Ѭ��_��`���B�ĸ��.q��Cy4�ݮB�µ�K�rn����sq��5����<����b�d[�V�M5�G0��䰴�0I�(��]��Y�fN�uJ���M�Q,&�6l��D��:��,�
Bj�l!f�g�%�$��%�aL�z)m#�̊�9��t�JNX6+{d��%+�s�SK�\:9�p�th4�.u1g�ANL-9��@�m��b�nM���1�B�
kɢ�������C�B���9r�Ԓ��y�XC6ռsf%��U㦖�!�	7����yqx\����3BO���Z���^�8r��f����H6Zߡ%w��D����M�Rr���XAj8���v�&ƅ0�u�����[w1�{4d�\��ކ��R��/��-�]�6��zI��#N)a�ͬՙY�w:?�
��I�VXJ6�B�4�ir�(r����MNef�ps�H�����p�yd����
2�W~�v�;�#�+�,H��i4֒+�ܶ�/j
y�lx\$1h�T�O�����M)�s�x�R�X^����97GWG�UX�v���Y�Ng���z׌�@��x�M������*���b��]8�wg�4�o��5sb��1n���@ނ� ���Vm�(d~�Y�u- �Wk����밻��q�Zκ�]bܸ��ȁ�@)'ƍpvɱrr�YKNn�_�K�k���f�h�T{�6��V3��Rmy1�Z���8%h��j�Q3Ic8��ZBf�r=D�g�f��i�jm��w�̔T�RK~ё)B���qp�Ե@S�9'�E��P�
k�y����R�1��X����u�,	0j�OMI�,r6rx����0Γ�ҥ/�]m2� �5��P�
��J����2�F�}X\C��ׯ��X�x�9s���R�fEW}�s��p[���̛b	[a-Qs�0�����*d�Y<�|9��H��w����
�kqN�նh�T�-���z�.YTûm�;�7�UXK�| ���u������s�L���\39�!5m��p.�����SJ�b�.9�?_tbÁ�°�1�d}�s�KĈ9QϢ�(#�lZ�K�M�T5r.�ɤ&-���l���]��3�9 �b�Wa)q�fTWs��b���r9�dE��Y����y<���o�K��/����H��Yt�{����)��ª�\�0r*�Ոx9�֝L)A�DN��a�V������Y߅����W0��E��r�V��w��*,��f��!��ڵ4W�4]�%�Mq�lĜ2p��.�-l�|q,�j�Ж߫.4dJə�f�}x�q#\�]r`Bs��d�5K��ٗ���9�n���ڒmf5�b{8�[�7�^�n*^�a�Z���a+�%'���_w2l��2���ME�	�6��Z�1SK�2�I6�7�<5f氹VU�KV��ͪŠ,l����R뽁��Vu`܈)<9"��li��SlB�7��؃ǚ-Pph05ѭX.k���%��"Pہ�
Rvyip�s�/7�jUk8��7-hw�+�_��H�B̉f�^��ōY��s�V�Y���f1f��n^�Rs��S�V�E]��_7)��YXK�t3�AO�Ͳ�s�K�M-Y�z�nx�bڍ�vA�!sa��%h:�A�M%����6@���Z��_ ���fʝ&�(����)%�r g�BӒ���p�j`L�i��q�ה��t3�{�2�*,%j��^-�.Y:j����˃M1O��sl�ϐv��Y��uu�7�U�N���Y�bάU\�c�Wa��_3�Xβ��pY�7��l~�)��Y:�\�ϋ�+�Ѿ���qS9����u�s�ֻ+�������p֒��qf�i���K�����U���G�1��[jr�lv�Js\��i�<֝L��Y^`�\H�vۤa+�%lޡ����Sr�/6K��	����,��M{�Z�r`��C�Q^Kج�c�@��-ц�ܼ�G��(ga�,�ͮ��#nٴd�� ��[j��%{Qּ�u�6	��3rjņ�v"˩z^��C�a+�3h�#����)�,;E��@1��,fs�~⪁�%�}���猚.Q3�|�uu��L��%�I'E�-|ɦ������}aI��h%b+����ΆM8�F(l[�!X��!�I��a,�Vr s�!sB�Y74d6Ba���݋��S'L�a`���`Ȩ���6�H��
�rȠY�p��YO2d��΢\�u\�8`Wa-�jE�p�Nk����Z�ž�|���͒��B͂���8�M�w/��\��t����M�fH�����j���}����Vf�-a7mK�в~KWM�Y�,0f�^�Z�^K̑�!0%��֬�F�Ԓ�2�n���Ԓ���^�jI7�VXKư��C�)�7����%)GN����۶i5%���� &8Px4�y>4��.9���µ�ĸ��Z�����jJ��9��l9%��l�5s�j�Z,f3�6՘Y59c��ɔT���Z�+�M��*,%ۜ�Ky�\�.���m�Ԓ�O���3u�k�[bf��%nVec�rِ�[���Ƣ�(�7�UXJаY.'�.8��M%�ґ#���>�a�2fæ����2�M��#sV����ؓ#��L�a*,%緛�����������b�s[�n�G)�%b&s��Z34+�0SK�[4d�r�y��*�%K��^!5��d;EŬ��4��� A�X�67pqȖ�+ܬ6gu��W���:��u!<�	{6$�Z����Y�뿾p�wY6bΚ5]�*��\��\J2b2CŬ�%`s��Ԓ'Z��M,��S�Y�fȹDf*$����&3X�̪k������V%O�V������DSR���u[�=6qJ������t4�.9kh����+Jl�殬��W���[nz��R�v`�ϗ��q�����đ)\��d��9��,��֒+ GͶ'w�C�y}F��SlZ�h,��R�f��F9��h�#f�V�h�q#\��D��sfɺYd�*���9D�!SJ����ʹ)D\����M���h�p
ѱxp^2q�
Wa-Y�g��E�첟R��M�D9<[����3�n�/�ؼy[7b�M��R��0I�(���D�I�1| �<&m�
#�,$�r#h�,=6H�������jԀ�S�����9d�<�"N�@mJ*H98k���}���q2-O9n���N�6z`ȨΆ)m\�K�l�𳵘c�A6���K�lS���6��n��9BؘYW3���G�3�9kŠY�H���٬�#jp؄!e���`sOo)2aJ�%b��1Cf+0=�Ѥhga˸��"�`6aJ��H�Cʰ
*R�h�e�ei�sWo"G��$Ɔ��:�f3�	�7��᪋T��W^M�ʧ�.��.��f��Dtb���4��D��Ԩ	�|a+�V��Xض���F΁|Av�f]Ò6���JQ�nh6��,1a,|	.��fk7b.�9p��^�d���AF���	��a,�V����ں��,"7h�6h6l�K��V8r�"s��,Ͱ��//ڣ�.+)���s���3������J�-"V���0�U`̸9����~�d[a����<l��V6�b����s�&<ca�����^�^8K#)c˺���� fw��ta*�\Ì0%#=#���7��/F�0aZ�u�%�=�����r��h6��;}��0`Ԭ(�Y15l�T�	�W�b���������ƺ�6EN��p��o9/�9a����ln;8n��0X����K)��eaD�0ܖ𤌫�hS�a+��q��y0n�(�1{d.42��Md��U�I��d��}#��%�f�#e|]$�0le��9˭�Aғ*T��RL�xFM�S0��d
�|�u`b ��Ȁɕb��a�����/;4�1�^�p��!#�`6��{��i���E.�4�X�f�I����6EN��pj�3筜�����f5�lMX�L��Oϰ�e�E������&��$@6��mC�0�W�8�����Q�	�|��Y���&&%K¦w8�.���s�^�KM���F�5r�0�W�,���kSD��?�?S�:0�l%W|P_��{.�8\��3n���g���������Us��0d�U�b�P�&[Y���/�p��w�L8��E�#	�VF=��|�7�.d�&k�X���fs��0X���>�K�~f�,����FLxR��E�)r°��S���q��0ʾz�V��a�G��DA�t	_��2����l�Dȸ��vDN��0�$�9��nh��Z�?.n̐���Mr��y	.l�,�E����T��ca�1n(6f��P�M���F�5r�0�W�����	���S�"�tp�&f%K¦{�Ҋ�Ė��-�$�<��mC�0�W��nj�݄Q�[�j^1j�<���fŔ�K����fa�,4��2aJW���i�X^Ͳ�����I*Lk"��9cl��u`J� f-�R�\s��x^�Ე��2l��8�f��9�Vn��5����Cfݗ�(i���E�8x���䰑���_]D�"'[Y8u�C����ɄQ�p���W08r�`m�"l��/�f�lha 1	���.�M���,�:�ɍ�(c�N�^~hԀYnĸ��Ltk���'l)�pY�p���C������E�)	�VN��܊@9 ���@��柩D�Rg.lnؔZ2`r��x~-�%'��a�2Z5g��g3^�c�%`��Y�+����F*Iӆ�0b��86��ܜ�r�$�$��mC�0�W�8��qg�v�&e���Jp��5b�aR�$|z�1-������l���q��m��6����,N�u���	��d6'f5���d�ȉnRLI��c�ĕ��?c7{��%m|aD[Ð6����,K�(�Z�gl�� ��T�L)S�V4׉��/.K[�7d�,P�8fI�9��a#fIP��ԝ����(i���E� �΂f5r�A�@�#e|]$�0le��9�p�A�{�&w���h�,|`Ĉ	��������j�l����27���E�)r°��S�8�ׇ�2d԰	����fՀq�f�D�H\E�t
cJ2�z�On̠A� ���E�)r°��S�`�f��9���A��\0\�,7n��R��m��%��ͽ�L��4m���Y`�����-�p2�,�m�Ӆ�,��ǡeS��FL��0r�I9`ܜ�b�[S.����,�M�����)mlaT[��cax5��rɳ1C��NI���f�����FMdS�a�1\��py��1�f��Q� ���Es>)�WF=�����EL�r���L%��d<�>0�x���xt/�\ܰ9��QF��%g��p!g�/2o�#�2��̢��f	��Y�$M�%f��Y9l6�@oڍ����/�hk҆�0��e��M�G���	�Z�كٲ��0δ���¹	9븡�Y��0�cax5��+�F�b>|�Y�dd��J�d|xӚ��?]�,Lb6�0���ӆ�0���]^1�Xtb���
t�&�e�%a1>�i٠�C�.����0��+�lk�a,�f!@�����l̐y[t��T���aL�xn�&7��� �0�S�Ш)�WV��<����I*Lk}0�������& `�7����L%���22���[�\)&��r�e��ټ�ͳ��y8U�/	���Mˆˆ͈Qs=7�����/�hk҆�0���+g�Ő���1c&�eq%a2>�iɸY5ׅI��0%���lcԔ��&! �Z��1h�j��D�$�"L��1�}>k6)�b!��MX��F�/i�XVm�.�&v�J���
g�:�%a2<�i�,N4n�c]���0��+�lk�a,�f! �6j%1�P�3j"[W&�Û�0�έ�_\�JW���i�X^Ͳ�����I*Lk"fF�0�Q�r����8�B5��D�R���B����Z2`r��x^��"�:�y9�������g����&�����Y�Q�1n�F̈�R��ca�1h܀QCf��)��q��m��6����,*��e���#���D�,�$LƇ1�2\�l�eG�ɴv�H�0���H���jny7pXg2`���.��1�16|��p�s� 猅sX	G���h��!e��©s��_�u�Cf���b\td�D�"�$<��7�XBn6�t�"8�IW���)�W^M�/�4rV7��#������U��а�D�掬�e(FN�R��E�+r��ՅU�,�"G�~yR�
�Z_BF�0�Q�r����8�B5��D�R�T��NL��#2p`0j6�i�GS%BI8�sZ3��R������XX��F�5i�X^�����3�k�&8�-�+	���LK���Y8݀���f��=
#���a,�fa�w��,&1�as�.�Ȗŕ����ɐ9]�,Lb6�0���ӆ�0���]^1kǍ9n����i7n"Z_�Ý�9d��np�,�0��+�lk�a,�f!@�����l̐c�Mt��T���aL�xn�0Kg�K�L�䋩�lhԔ���YE�H��
��>
I�TGM�E0��d
�|�u`J�J=-����h.�W5\���Y �ȑ#�����=����q9M�%�f�E�E�3n���i�X�D�ͩYڛS#F�0��+�lk�a,�fQ�-�}0�\9����Ȗŕ���0���y5�X�4p�p�.i#F�5i�X^��-��2�x9�E6:� <Ɔ/.K�̲�s����p$���fKR��.�:�[�Y8d��Y	5o"#&��%�14�i��2t��b�I8�IW���)�W^M�/�4rV7�K��E�$�"<��5%�m�̏f	�	Sʸ��vEN�����Q��/O�PaZ�K�H�:jZ.�����'S��3��S�V����V�R|N�r1��.�5kg���L4�+�!AXS���f���{��3)���������������F�4�[dp�ZW#Ø���YfpȰA#f���u��
C��ՅU�p˳���#�oN4A1�"<F�5%�%�I7g�1jĄ'e\]T�"�_]X��<h�ڍ2b6�)5l��fE|E8�sJ5h�l
�-�]�IWծ�)�WV��O�-���8k����)m×n	��)1l6�f��B�ز�EM��pꘕU��/O�PaZ�Gf$	S5-OM@�lo��)T��:S�j0�L�%&W���.�zA0�f��Y�nȬ��A*�����Ȱa�
6\�,y5j6����P��_]ĊMl�P��2�Dx��F�/i�XVm�b2Z����.�5AFMd��J�dxx�n��[cfhW���F�5r�0�W��W����F�Ȗŕ���p�=�A��nn�NX��F�5i�X^��.YQ7k���ac&*u�K�d|xӂ�C����n����E�1j��ՅW��o�mj��٘��&�5q%a28�i��Yxżh�p܄+m\ad[#�cax5��*rD�#I�0gk�N�7"�2���\��hG�
2�[m3d���N�ͭߘ3p��A��7�g!_G d6�T̬�4�]:��|O��L�h޳�� ���,�uYRW+�K���U蠓m��<��W��r�������ŕ�������RBCf%n�7l�fn���pY�wc�����������Rd��b��Y����*2�·^��Ԏ�K������5��¶͠	�C�n�u_p^&���,��Z��6�C�n!�fI�/�måU�2E�H��Γ*T�\1[0�����0IҴ��d
�|�u`J�R��s���
�v�hUɈ���~��n̬��K������R_x� ���� ̐�R�ӆ�0b�.�Af�p�
5guX��F�5z�p�W��"Pa�w��,��Ds�C��jY\I��gZ4\jΥ�̡#,i�#�=m8ëY8�ݰ�UDcf��t<0lĬ
9��f�d�ɬ���p"���%f�,�%���­&V���E�1r�0օW��˷	9���7�Y1Q��/	���N��1g����0��+�lkԴ�,�f! �J�#G�2`����Ǖ�����ܘ6�e9aJW�֨i�Y^��./.�ic���M�a#&�e�%a1>�iɰA#�9b�lK&\i�
#�5m8ëY�W�#R�Ii=ٸq�f=Ռ�m�9�����Z�Y�f��-O3dn��.��8��,���M��ag�,�峠�Ǜ%�f�b�����o�{�[.�e����6��ˊ/�܆L��|S}����la[?4!Q�����V\���x��P|�Bsk��*�	��a�"�f�����I�0�I-��YT��Ǆ��{��z?fo �����mN�@ 7���Yҿp����pi��kMfف�.��]%g���B�Y8j¤Q8ʂ.}��,����M�Lw�2]�uX�`b-��˂/�ޚ���Չ�{����Y,�@s"&�G�)G�@m�H&L�uPA��$N���\�\ƫ�Fn*�V��e��7jܬ�ʝ�j��3�Jr�pF+ټ�{��0G���h6FOƺ�j���8!>�V��r*�ʑsp�hI\ExcJ6\�,���0Ǹ�p����fW��a����g�p-堙T+6B�frf,V�V��²h"T���hj6���%����G���hvEOƺ��ny�pQ��̈9��ɴ��"�"F�9�0l�2���lr�'e\]T���c]X��<f�x�Ԍ8�Y�i_#ÜR��E���g�	Sʸ��vEMƺ��ny�,��+v���
�
�q၊0�D��ň���r����-�,*m#�_YX���+rD�'U�0��-I�TGM�[0��d
�|�u`Jي�1�\�څ9W���7K�҇G�H��_�M,�%;�Y1`̼d��Z�%(��6K0JI�6��K�ͪ��Z���&	a,�hk҆�0��EDG�xnȈ!�V+��%�Ȗŕ���p��ĆN14`��)'&,i�#���a,�f�����|tæ�lȰ9D��ܠY��ب2�J�Sa�3\Ȭ���x�Y�D�Y��0�cax5��b���~m��9���j||IX�wZ5?��1sz���&Li�
#�9mëYȻ��������FNt��J�d|x�n-��9�����0��+�lk�a,�fa����Ш�p�L[D��K�b|�Ӓa����"g��ȁ��q��m��6����,˫��_�T���L[0�������& `�7����L%����UQS�Ȁɕb����uaF�]w#f���E���
4[n#�������]<n"��H��h%p�l��SW8K+)cˢ�=]��«{ttD�u�c�9f���j{LAx�
_:6\%�CƲ �MN8��E�%)�WN�à�S�Q���C6��fe����[�"/4Ss�Y���5*bS]�
5�w�,37�)ƌ�8���.�]aH����ny�*������h����è��:�䐑��3`��?LuQ���2|ua�3�ʚ�ǌ8�fK2pЈ�H���p��4�T�N�R��E�+r��ՅU�pˣf�������4lV�
�
q��0�����,s0l6�t�;<Ċ��J��)�WV��<����I*Lϳ#I��i�hf{C�L���T�L)[X�}8`J����b��z�Ásw�Y{7j̬�g�F�5KI������0�8d���ţFL��4m#�,��A��M.�e�NX��F�5i�X^͢�-Z<7b����̢�ٲ��0δh��YDjN9Ko����mC�0�W�pȫF�0rV�̺w��Z�oP��
�ƳY��f���Tg|�
#�,�%�D��Y�jbeO]D��_]x5	�|b��q��r̸A�1Q��/	���N�y0b�:8C/3aJW���i�X^�B@ޕR��M��|�D7>�$LƇ7-��� 2n��ٓ��q��m��6����,���"G1pf^al�D�,�$,Ƈ;-��ˁ#f�ٖL���F�5r�0�W�,�"G�~yR�
�3m�H�:jZ������'S��3��S�Vr�$Cf�(�d��r1�x�f��9����f��pYlk���,7nԸ�j���H��ކ&JI�d�*�Vg~1jp7Ca6�H_��0�_]x5	Z㣑���b��9j�D�$�"<��1%�S~j�0äp����fWR��.���C��[m3���5BX,l.��
7`����R4*�O]�
5\�lf	�Y�ۢ����u��
C��ՅU�p˃f1�cF�4b��ɴ��"�"F�9��l��9iԸ!��LxR��E�+r��ՅU�p����Ԍ8d	�������aNy�ބ��S�?L)���9e��ª��Q���Ձ��"�6�*�aL�f��s����͆�h1eQi5]��ªoV^�#R�I	�˽��懘�6����!#�1hf�m����ok4�Ac�1�|�������B�΋� ��y8���f5�,E1+�e���&� B؄��8o��v�|���պ�����Vl��S�YT[�׶������.΅M��uݖ- l�-��5r��D��x�SM_Y7\����7�rrv3W�֠�fٺa�|�W�妸�e��ٗ�9fz�l����Y���5r��Bd�DK���G���D�[j+-禮��Zf���:�/Z}uwo�,).�M��2D�RM��u�r֋Y�bK2jRI�p9�ĘYX��4@��of�V���e�kE5��GLҵ�[�\�I]�;u5����̀Q�EM,'��RPᤜ�x�LV(11J���+TN�8VL�vU�V�d�H.bF8jԸY�p}�.fԬ���!3�Y���K���9���j#hĠ��l��A���_38\��7XC���w�/B6`Ԭ7����5
��$7+gcn�,��r�b%��J�Y�k�(H7kt���Z����Eͅ��h�9�����YnB�h�KA1bЬ豹|�Y�a�6h�j�ՈY�R�F]���>�C@��k��6̆�c:tj.�9�A�&�\E.�����z��f��x�{7���%�d�25j�p̬�r��@�,a0�_:�fsH3�p��bK=
���Ij��f���+�����J��7`�,�R]0n�Tb\�Tj̄�E4�c�P���ff�Ɨ��
ͦ,0p�,�]�R��^�%'g#	Gݠ�J�!/Q�)8fԀ�2v������4���b��p.ϊ��YI4d�)�fg�{�q��V ��˾LݬF��1��]�F�������9����� o��2d�$=ρh9�O�]8`�k����|���7yZ�5DN�0laf��fɼc<��"vn�UG�5K�X[)72��*z0Z4w�',S�H�ڎ�$L�6�v�i�/PA� m�I'E-횯�%]&vs��p!��Qs�^��l=ќ �-gX�.f"��i�X��l%��Kl�UÑ2�,�m�Ӆ�,����"N��$w%��nܐI�����9�8�Cƍ�b��i&�2�"N���E�X��l�[3fȈ	O��¨�EO�°j��P����VwI�	>ݬ:���u4#G�8�h_J�5������ԀY���p����fWR��.�������fC���j�+6b��ג�C���p�%�)�pa��4oR7r2�.�]aH����'���͒g><���
�$�͑��Md��U���aLif�؜�hĈ9��O�u��
C��ՅU�XI��9fV#|�Z�l����MȉH���pP6�)��Y�`N7�&,����jW������%f��$q��+)��-.�5 BF��FF���L�Z������=�D*YeB�hI
oa�,�3氬f�.��%��w���p����-ȰY35j̨�%���Ѭ��0�.Y+4l�I7'I�a+�sw�cFΈ5%[-99���U+����F��S+Đ1����Z��BfS���s�f�,���MN��p�u��]J7t�t��sn�r�`���R��d�����:s�s΃����ņL.!3ebn�.yn4+����>\u��̹��+&f*�l��os~_�b˕^�bĬ�7]�`.�Uی4K������4h�d-�4���S L����F�P���<G��ᰑæ��-�Ų��t�q���`'۴Řasư9�׀c��=zY�UXQ�5Gמ�&�z>�2ZxFK�jp8�;b�H3-D6#�ɳǦ�(<'�Z-��gf�ՄD��TI����mu6Ʀ�.XK�lnL%���\���9�+�:�Y��P9���sW͕0SK.p0r��usc�yq���?7I�VXyA�լ��J�p�,6�;����� �k�M{6���G*��h��[�]+�9Ԭ�ǂ;�*�%�vA:�nRM��@��⑳�N��KBfۅ�2Z,]1p�߼8�\�oS�8�<fڶC#�P�,W�Mg�VXK�\ϫ G��!4wx=o�|��d�Eγ,�5Yd+�B<k��<��t��������T��Ȝ��
K�N�č�;�|�7�����f87��
1r6�,\/5]��]��`���6p̼{]6˦ �Ѿ��5�D��j�����9Zȴw�2j��K�.���KlCe)oTN.8 m���in`˅h���L��a+LK6��#����Ϊ�N�Im��z�7]p��,���(��z5�W�V�Okw��<Y���)�|��[o�<�з��<tl���
g1�t"3'�
s$��&ӌ�7w�pީ6��yf��ϱ�Oa��A���kr�亙���s�Aj��'ޒ��%l_�fA%S*.��y��^�Zp�N,���� �髆͡�۔��z^L9n�84]Bf)l}x\���S�9�/��T�Q�!9l��Y#2m���Q�\�{�L���
3[җ�F����8�ޙ岜����tg�*�qSK��U#s�"�K�~�����˭��f-Σ�0FN�a+�%rĜ+l��Z�4�p������u���
��&V�p^�AC$9�7QJ�&I����%p�,f2�8���LX҆�0b	�M�Qc�%��c&,i��� ���-7�&ZZE���� T��xj��9 ����؈�,�C��u�'Li�
�䔓���l�0?,i�V����k}��1���JW�%d^��E���,<i�V�D1�r���n�ᰤ�/�hkX҆�0r	3gցV��C~���V[��荙C��Z҆�0rId�c�K�py�Vo������m#��l�X^H�[B�hIz&3\ج纮Ԃg;8팚S{w9l��D6l��Y�'c�%�s��V7bΦ.qsؿ�p�LM�������LI����X���E�e.��*/ׅNMҍ�v��^�fؐyl3�&9�O�u��M-Y:��%%��t�,�K�fj�t��+'�s���d�,�5gcF�2N���Z�F��|ٹ�n]"���!#G�e7�py^7v��KJL)��rVa��N-���
[ Ϟj��Ɗ=%5ۤn���K��rE�ѥ#�2���^J�da5�%d�Y�n�"�&ZѭVb#�B�g=V�*�T�n���y}��I���Zr�E�񬭬[�[.��~]��U=2�5S���[>�&��.Y�lxq�9F6�%�9OU7[$���.��]�pV�ү6-���,[9�dm7bܬ1S�x�̅z�j�'G3�;&w����� �n�����=6몦5X��Yfn�u���Y���Q��ݬ� ���XC5U��wp[ۅ��i��[�y$0r����.��`.�p�l�lZ�S�P�55K�*r��\8���H����%sA�=+�fM��Nv�u��|��jb8��ZpĀ9��5��b�s��f��%'�g���� �誊Y6%�;�l�\W�.Y�[��[���>\��d+2+|)�C9Sg�¹hk��Y�ݙ�t�OM���O�hOG4E�7�1sgVǍ�)�06���&��᪫�/E0G���+Ĝj�bc�X��^�98/66`�L����j�Y��CLM�6{p�䙊fJ�<��.�M��S"l��d����03(��͡��Su��h6v�E�n�7K�8;��V7�,щ�FN�6%k��%Z�hb�[a�l}�W�����.s�m��BS�X*wBͺ�Yc2�H2�ʟ=�	�*��hт������{r���t#l��dA|��G��|�9��5�6���R�t]��oڑ���.�#jd]��h�pVsb -l�]��+p~,�s����U�xٯN)!sd�9���S+��݋�"��5�d��b�=h��@pP���a+�%�Y���f�t�\J�Zޥ�G�7s�;��o��dEn�R>��l5�d�p�\��SLc3�N�%�F��eF�
x_v���\��5�Zqr�9�]6U6�ɜ��W�Y0؜�p��&Z��`���.�����Y ϾCa���f �4d�Ԋ˰���2��b�A�LC�z���fS�jU2��9�.��Q�I'E�-�%��9�_���h	nf(s�$�W]�X���^rд��kf˫2¯6n����jll�.YK47n[1�Z���\�p΃j�:,`w�i'�0�UVV��E{h4]������������36��#f
~����V�C�9n��l��p֒%�����Rsx��,ڃ��Zr( ��l�cku�։Mc��bf�P�%f�Ԓ����\�1���Z��,����<H��z�aæKVc��_¥WJ����ALL-Y��/��ސ2U�c{�W̍�E�t#l�]r��HV�7�Hdܬ�5Y���nz��f��L��uz��y��.��p�Y12�O����ur�n����,s6+����T����b��Z�K\ΧU'ӈ�s�Ь���$�&��A���P�6�~7Ǧ�E��M��X�K^ �����.Yn�|N�	�Ԧ�Uj�.ۭ��<Ț����R̂:03��6畜]7��8e�TXygh%��C��)�r�ߢ#FL�:�z�Y���D[gjVe]Y!��-8���Z�����]�$K�0֒Sd��ש���G��5�s��f݊=�Ԧ��;UJ6{a�9ܸ��=���n�Đ+\uȮ��e@F͡�+�<�s�aS+�\�53s0=�v"5g�AW���K���s]o��Z��АY�Ԑ9�Ťއ���\'6�+�L-as�ai-YěDs^0Eh[,%7�ۆ�t��L�fW��ʪ�ZQ9�s�I���Z���epb��n�9���3��.9�7wv5j*>�q8bF�'�%�7[�9��T,����}8Yr�$qR���%j���+df@F'D��%��H2k�����,��c7bМ�
��F��>�01��nf����X��̐�%h�노n�+�K���j�%�i�.w4�^\k�fJ�\��%�l��I���Z"g�뵴n�g`�yȬ�9]r�^�S����%���n���&Q���f�~�K��	r8^ �$�[aZr��1|�G�6G�i|]�V2�2d�c��"dܬ�%bS+.��Y�7�P��W$,�)/��ܙ�V%��er��6)�<�g�#�"��0�8��Lk3�#Z��Zr�O��ǱdOa-9`�D�b1S�f�\0��3U�ŴN�u_�j�z�96�H�R����,@l�L)��f�Z>r�n���KV� �ܘSJЬ/���N�	��v2�h�76��2�T���r�;3%�u���/61d[a-9T�y\6w�7�Py�=8]B����`,����E(�d�����p�>�Y�������!�Sa+�%GѢY��_@
�6��a��`�O���b���4�D5fҒ���6u#+t���eF&ƍp&J���f��߶@�سt�\V3lj�:�9(�N8��znKfs��A�Y���k�lN�"a)̼�����pJܰ��sݨɬ[ۅ�(\z]af��;i�2�������Z�.9?�p�ag�V�b��6p��9U���:���[�e�"t�\4�sVw���0s8/��g��<�1��l^Κ�1�H�
S \nf���������P�"r}��6,�b
g�3gۚ����`�I���M8d�	H������qTtE�y#���z��.0�ܕ�@��U_�W�1��]�[�FM#j嗖6�mؘ���z�9�O1]�~�$����$�[a-A#΂:;���Ml�`�DC4nj����LZ�p�4��{W}���p����fQ�i�G���t`�Q;\u]1l^�w�]�7�c�@MfMĠASK��ݍ�qSK��MB�ȩ��RΑ��b�S��h�7S&����-�,1g���P�,�C��s��Jۥ��M�9������E!�c�/�d\j�88��X����Vpڒ̀��/��7��|���(Y!c��-0��VbpuFF̨)0��GТX��%g��6��0֒ͭ�ws���b��@�����u M�Y��������f�[ ��I��\8���O���.���#��D�cM��!�rE�F��.�7pEN�� rI,�T�Ɂ���b��Yq4l2�ݸ�ԣ���P�
_b�ˡ� t.C3j2f̰�#���.sm� �^9n7nj���B斮74�ݬĚ��ɤn���KȘy䥾���-�{�Ǧ�̆�^�n-1����V�.͙�<����o���ےY6I7�VXK���������lg���q7E3��s�V3S���Wsd-���f@�zml�c*���>oq�"a+�%�T�β0s��r=�.ې�����;��\�`����~5#h�%G�d��.� ���/h5qn��0Q��]~p�L	6���_�:�i5�_2��W�9?��[d&�S�	z&֒��.�s�1Ù�fܙ��63b���A���IY�f.�V�@3�<2)��z��@��O����^�E�V�1����$�K6r@[J�F��guϾu�7%[��Z��[��&�N�m���{=N�X�OaB3l���P�%�f�ɼ���`V��·i0�r
�|��n!g#g8C����}�ח�q͎��P�f����Lk���ʕqs~uɲ�s���f@�K��p�8��9e�����%ې銗��Ⲟ�Sq�~�b�^8�.���Kn��m�rX�����f�w�����f���50W�KЬ0G�Ȱ�%g�M���\��d����t#l�]�`��<'Y)q3SU��Bv�]U2٦3�� ���ޙ��USt��N���P�
���,�S��)�8�����R��[�b�u�[��z�Vɖ��^��"ϴ^7��f�/4I7�V�1\6Gf`���˘Z���eaF��Z�>��ɵf��$Y��x` �p��¸�ݶ5BSa|Y?�����a,��7��wn����&�YN�ʺ�Ö̦���BT���w���b�O�f#d&h��گ�fVdY�?I7�V�%lN0�t��{��լ�!~aX�U�{;�53���˴�Ų&�n�9�М��Pө�G�v�w��I@j��}N����wJ�t�5Y6j�dG�����nڴ��ȜY�\q�-܇2Ͳ���.�e,&��0�%Wls��v�O�u;R�n�0�w5fm[s9��l.L8ō�y��,\��)Y�f��o~A[2�8!�(A� �._����k��dj�W��j���b�K�n��Z�9�K�,4���c��t�by43g��খ���9�{�����/gY��=��a+쒳|9b����K�ə���갩%�[;0��a�M�\0k�po��%y���iϦS�y5�]0��a+�%d�#�C� �KN�M��j��)d�b9Kz��3��i�&p��IK_�B�L�ܦ}�lj�ĸ�´D8Gǂ�.�y��"A3��,�Ó1�C��ͯ���\2f��'�Jn7�@�y��VAL��*̼��Rޘ7����r�CX��V7i��d�Wr��q�&�x%���Wæ�\�pN36��z��%Wx
3�5+l]ŌA�i-��+Ő�E3�s���%Kl��E{r"BC|ɒ�$����v����C߶aJ��h� ���4޶H���Uc�&sR�1��D?���q��qu�����r=�N&[�z.�����6�p�ga� 9j�,'7��K�,C9�˰6I\���V|$�f�֌1��Asٜf*��9d�٬־�.9p����i[���9:.�
���گΊ.j5مp֒K� ^o1r�T{��G6�"�.ٔ�{�
o4ө�Z���u���Z��ݬ5��JզC�7bT��I�!���d�,HǓ3���*��o!��,�5d3�VN�ȹ��`Đ)%�k�E��Wa�����Zf'�}�q#\��dYoIf;1_�4,o~=�Y�eĦش�tѠYe0w�%k���,�KMʩ����Kͺ�_�-\���ʉ�T�
k�Axi�9�;8�n� ��[ݧZ�/,f��@��lcs�R���f�fc�%a��5��8���K���VC��,�vcC�'�1ō���o��<��Γ���'Luc���YḉT�A*��/��x��C�,r�0F,��p��KȰ9ẅ́%m|a��fQ�c���0(��T'D��%�m=��G�Vb6�Iͅ��`�����%��xt�C�6��I���/ؖ4aI���%q��)mx��OM^7\�C̶KbE��L�<�Xr�]�{��q�]��nJ��33aJ�%����
Z�b�,P��	���0bItxgaxy�5l��1Fκ��'6��)bI�ca��Yķnq��hxd_]��0����jU>5kr03#F�J�3�E+9�����Rx<B�hI
oa�7��#�̲Z�u.%���'s��M�s3�� �������U���!3�F�Up�B�
K	�%�fl6�+�3Ch7�4`��Y�r�6�%k���s�/.2����_4�T�F͍Z��t!l���*߱Ò��]��`k8�hur�3�^F{h�47����
ݮ��Y����]���Z�}!7���[�K��x7�wϺD�J�6��]���rr��ܬ@9aJ�%a �0V[/�3d.Ux� ���KĠYo5`�Y1pȤ�ca�1�[��uasT��%k+�3l��'�Cɂ��c��dJ����;쒵��G��^�87�TXKԜlԐ�,�.����ac�M)8v�,�AYC���h�^.N5OWJV�]]W1ME9�q5��}!��>\���̕GsȘi(�΋f�Z�3E����<�a���́� ���R�7c'��0���o8	�caC���f��LI���.�sQ��]2�J�%a��0V[GXbΌG��V'D��%�4.̽��圾�iu�\J7d�0p^bfŷFsV�'JI�6���K�lq�.�ӐM�����poQjV�!,i�X��@sX_&`��Y�p؄%m|aD[Ð6���K6}��Q�����q���g�9 9r��	K�0F.�?a,l[�\�nߍ5k��a,�X�cad8��6��ᅴX�%����gZ��^4h�H�ɴ`.�g<�6
���q��FM[�F1�p�޲�n�,3��K���~�Wb��3�d}WU�R[#8��|��Y��,S11އ��V,q6�[�T7��m^4��̆�Rq��5������bk�blJ��W�Z.*6rj(97~!Y爙��UXJV��d)�iB��y$���flȔ�;����Y�U�ջ��S4r��� �ٸ��MW<֢4��W}�R����T̜�d��K���ҿ�(0�������c��N��w�����T��a�b���[�S��b`�ʼ�`��5q^����\ɥ��:n�Lʢ���)[*<�ޥ��p��\6Ŭ�m}W{�z�L�v}�r71.����,����٨�1���--4�d�Wc�Os9jR�\!j.V�X�v=�Y6� :�q�*�%`�w�˱Ϧ�X��%s���%�6\�]��~�ź���0�[a��y4�cFM��9����'��������a�VY�n�i1�ϱɬ<�8��U�%㠘�����᪫h6g}�d0Ո8c����%�z�
yթ�FNX҆�����C���x8`�Tƹ��*�sd��&\i�V�%����6yiä|�
�K�UV�	��@	B�'L��1}��8`�l�`�N��S{Vi�x�9ȯ83k��?����u��~�w9�k�+f/z]��i�F�L�m䬊����jV0�C�k�TGf��\�헌�׉�ul�,���ù�v9�Y&��+GL�N�
s�YY4j"���,���=$��_�d6~[��9«�k	G�R��������"�.����f��y�]2lB�.:�#�-4KK��f�Z��d䨹f�"j̒�R
4k��1urVa%~-76h��z��rV�&�;�V~Ymr0ퟘ�n��`�$ewF�;W館𿠭��`Y���u�d�\��ֹA����:���3�q]�z���]�币�4dVaA��+r�Ѻ��9k�L����/�",E��: B�'L��,1}4`_92�� sڬe�Yͫf�լ�3S�ތ�먦���������(uÉ�m��1Y�x������	������F7��]���L��E��u���n��ep؄H]4����T
)>=������@���d�e�I4b2��4�3Hxd3���:2�+x���uz3jN0d�sP�A-bݪ-���f�\75h�E���s8v��L"}�L0��ڬۑ���`|����R|��25j|ɳ���B�R��C�s�6h��G��lx���Gp=��br�*���jo�F������r���Rgf�,Q6�vI�����as0 ���-���.�ӫI�k!Xs8+gm�TN��B��,�n��4\�ʯ��쮴��m�E7��BrC������I*���j6fTK֝�n�2�����.mAZ�Evo��q���q�]�o��Ȅ���^���Z!j��r�]�nbH�VV���1���ߨ54���΅�zw�L���s���s�KYtVG)[�Ep��#7IGq�0���J��`6h��_r�Ly�75l^s7t�u�c���ù��4�6'�m���/hh�w�����SY�!0aJiɜ�?6f���z��5`A�M���Mޮ|5����b��s�&�)
=�:�Y8)4)��v�����&Y@*P�8vW���V[����t���y���d�af&0.��dظY[9gD��̡o/1H�s��po�͠1sj�	O����pF�
������"A�׭��m��.[�ȌA�'	�/3#F�%^r
nՈ���z�����g�V�\\����V��[O8T�/S�f��9��Uv�Y��7�0��f	�YH�	6a�h���h6l�M$u�d�CnV����һ���B�FM��nV���f(�d\�����I�-���nh��Lx�6g�yI�������z/����n@w�^�
�bܸ1�1`�M��nΧer��a���K��3���[�?�C�ݜ?�������k��G�6e���:1����`J���{�l�]���"'�f`�{ʬ��]���m�8�^�reSq#�����;a�ט̕亩ukq�7�A?���kpVNĺl|�b�R�lb�g��fFM���.:n�(��ٺ?35ᨻ�hN�uC3�.&b]����s����s.1lb�6�khf��T��p3ү-��$�cs:�!��ps�͂�99+��j���ܪ�b��M���p���U�bd�'�u6C���Q��w0��@c&I�������
��q�Cs�I��Mk�TWJM[&�,<�1s+����j6tR�O�.��-lKkP����1��L���D����r5l��-��/Z ��r@�fC��bacf�r�F��N�SA�ջ0�,��S#f*��&I�K{Jx��"�@]T��p��f�^�k'MT�	C]t���u����,��r�z!P��Ć�5h6��+6Q1	&z]t������ͪ�	������f�O�?Y����u]��^��*uh�2�,�W�I�|�6���1}��H�&6�ک��FM����3hsb�#&���f)-+0'�S�H]���~!G�e���pm��7x3b��U��ə]�����[��3Cfl^�%�K&Y����e�����L�u��0/�S'�ֽ��ͬ�u�ڮĺ��g��d����[וb����l׋��nHX���"��Ŵ�~m*_��]2h>m0Lur�,��iy-�l�_����0�UN�����>�)����v#'�~TZ�6};��ޮC�!�C��dz8�y�����_:����Rf�|>%�W�x�ؠ���M"9�q��\4rڲw��P�RҲ(ug�z�-p�,^8	ߢԝ��j���M�UG��8���i����ޅ������
�gO�N5y����#��a��t���_�u_�K�� ה]�?��S�_�l���mt���Ű��Y��o��&�,�5]whX�Wi�(�uG��-6�g�o~��\ˤ�|�G���,i4]�L�
�l���d�����yq���X�Ucs�m��
��=�!I���~��WE̖��lK9��̵�TV�5)�#�]x�x��ܦDz8�^^���W�]�%m�^(�$!�a���9 �i��l��+�k''����g����G�ֱ��z��g�᜙C���MM�f=�u;��t�pΈ�<Eי9��&��dգԉy����('�[����E�.b�����R/hr�[dp@wx�^�&E��k�/�uUcf��D�+`f����K�F���ɗ���R]����fG�hj�"N�@mJ*H�<a�d�b�x���3�ڭn9�g�K��:����ưAs}��O��0�rY�&5M0��
6#͙(&Yw-��̉q�H]4��#&�Z&#벝>9�1�����vfc&<6/{72b��dвu�,�.�ph��Wm�M�1���۵_���a�\�<���N�S`��l��-��r�oli�ASw�-�e��
�j��̀�Fb����.�pԡᲨؐ1sz��ýb�FbR�_�TW�"��ZL�g�~�ån��͸)���LQkM��
?d�I�Z�5&s��8T�	��}�V�^�+�
d�S���n���R�P �#�Q����eװo� �W7� 2pn��mt� ��V͌���[0����Z���5Ur�8�bV�9�Ok�96癛$���er��庼ڿsk%�ueuk��V��#C�Y�N�fx��ej%E^����W/�ձ���I�M��[BOz��!a�nU�32�9j��'&��F����Rv�&:����%&L���W3���	���j��ʟ7պ���!��op�Q���,��oaS#f�V�43#̀}���M������u����ƍ�P���-���b�9���"oc7g�f�,��T\�T'��Y��C�b�.��7��Y�����KY̡	N�:1���G�2g3�]w4[�3B]�Aa�3s8?�lp�u����!��S0��jF�m�<su���́qk1I�݀qs�� ��D���-��x���hC�.��$���2=�T��n�/�����uf.��]I8rEɺ�W��IfY�!���説�CKĺ��G��nN1��7�73�W��;�)5�DNҺ(u���`i��B����3��vh�DT/�E0>��Q 	MhA��.��a4jܜ(�!'R]8`v�lt����uQ��b�+C� 8+�Y�^�A3 ݠ(u�m^�5;ğ�����[�%��i���T X�KL�:��Z����b٪99�4�uy��<2�nu��V^M�5�r�������!b��M.�ϋӌ����[g��¹q���P(��Ԭ!2G�e��27+�����r8ĴE`ЈY6�r;6r���!�8\��Z���l��u����)[ݻ{b��n=Oy9{kj&��u�Wsw向�&@Q�8!�y1Ks�ˉͰ%L���[�hV���o��-�����ܐ0pB�(*C�>�\n8����2RYT_���-@9��c3rB�.�%�&��ج?�~5#�L�t�,ǅ��#��/Z]tmѠY~n���!Qw@�I2n�]�n�Twr��d�M��(|��u�(4�j��b�"�}XW���?���������g���l�n� L�Ǧ���'�����02j������G��.�5_�5��A9|��Eg}��߫����B�M�:0r�ц����S�ۜ5A�Ń����Qm� s�2��ʣQ��O�fV~��Ynrȴ4���F��Dz2�f/�u����w�]���^,�#�eұY��f�H��	O���A���˹ml��>��܈��6�x��x6/Y1d6�bf��`N�ENm0�>��Y�sk	�+��\*H�<a���d6�G ��b�\�K��ȩ=n�<���ƌ���mf��17�RY>ۢi�`F���&�)Z��k��G��?Y�������%f]�
�|?b��RF��t�f�k>�QC��Es&m���Ss�l�H��nx F�8rN����A�\���:1�?9tv���m*�ݬ09l�:7� �~|]t �j�ʏƳJNx��,�M`nmĪb�"7���m���UKp�ŸY���	O�9�p? n<��Hud�X��rbX���R��_�6z�7m��m������C��qk�u���a�溊����Y����a-���p�$7��(�Z�Ew�̇
G]��D��*�\�mbA~�
_18����c3j�4nȔ22fЬ!9��M��T�l�4	���fM�44�Kk7pz�/J71ub�ڋx�VY�s񆈉Q�Ps�Yɰ�-!2.7����́`c�?5\��iu��)���n�b�ep��!�U�#'*��`��K�\]f]��f��N5f�n�9����	SY��*&����9r��!"�L�����9W��48wĤ�ݪ�_���7�&<u�3��a�m]٠9���+"��n�{D�Y�݀i�ϓSl=�aSI�Ĝ�Ky�`��!�:3����D��'���c$	��@	B�@=���
�`NR5�u��U9���$G��^��sN�P3o��mj�pL�G�j����p��9����n��Po����:1fȘ���I�E�-�LL8���,�9M�4R��W���Z�r��.p�qף�)�T̸	9>��r�/﷞��h9��f���7�d&9Z�-�mɸY�%I&Q���eifY�ƲS��0�~8���:3�;5k��E^ӯp0����Ĕ]��t%�J�li�Q�fwi�Ԅ�n�ذs�V�L��HudVb�Y움#&��+���~�jn/�e�l`8ɺ�|sZ-'4]wj�9(�(�K����#�)�u�͉�r4�Dz4н]~�ULM�J8�ly�I�=�o���lq�!S�'��3�a4���f���TN��r^�'�%�L~ܙy~7��+����&F54/3�hj�������W���ky�9�T���~5�ʦ��Xv��7t�Ʉ[��<�qS҇���	�����_�s��f�a��L�M�͍-6!sx\~�R��hN[0��A�M���$��0��u;I�k�B���K�Z�D�7�9��<AԲ�z!XNW�áQ���p��>8gF���Bf	��UG�:6C����uV�.˼�Vr����Ժ[0�}zѬ��cl�l�d=՜f��=|]�[l���f������+�ML"աY�+L�A���F�;�6s�]flb�dဳ7�����u�*����q}��0���D��p�9J�"N�@mJ*H�<a��|�0G�ªfP���3lj�M�T��jb��7S�9K�,2�SNugs�5sc��Z�I�f��4l�C��޻9�/�b�$�=���"%&�c�e����e���,Z��t�oMvm��l��6s��!Sq������I��l}7 f��1�+b�|���?j���[g3��r���c͗O��׹9���^�n"�e���nn�:�!��r6�TG0hJ݂tr/�{('%���m�f��Z�Ɔ�Z���ѝL?.�y�����?��fɑI����^bz�6�:�ꚉ3|��P���6¿uϗ��g�&�L����&��af��Y�aI�ፓ���΍��4�{�Vx��ȨY��>n7�"/Z���\}3n�i�L���_ʫ���Ve]�6Kh�,s3I�W�̈́�x��f�<�2Us�cH�<O'6�=1��R��
���>6aI-皸��NKE����ߴ�;�(Rw4�����Z4h]���ʦ1a�[FW�Z$ 6Jݕ�Բ;|,���/6hȜ�j��b��c0�M��Cg���A�,S��ҥ��M�R߬�M}�Vg͇��+�7������dZ(pn��YQ5���.��l̐�SH��e}�T��u���-��[L*�[v��e�*�T��V�B8Q�TZtl��P�,�t0}�J�ń'�r�g�Ѩ���ڋ!so^�:6wt�`#�H��o���Fs@>츉a��ʎT0`��/�Ø�e2��l��3�_r6<ɗ�.��đ�0�f���L�S�	��@	B�'L���y[`�z0�G�����f%kӊ�A��X�s�ײG�NK9�Yv۵k�|9o�����LR�e(�a��3\uj���ݲeR�p���SǍ��A���|��,���*_�ל̣'�6����u�����z����뺨97�|Z��n��M�Ib~��!p����x0߭;��&Lu����[	9n��E�[�|�nM�w�w��x>u�^�t�nb�ଧ3��Nĺ쟜袾�����&�����^�����;0%���A[�:��u�i�9Ne41�^36���T� 53߶�jn��o��5����ʈ9,�I"�<v3����3uS4n6�ݢ���]<�ۊ��u�΅�f�$Ab�����L��,�Z����s�ԛ>���e�(�ˏ{X�#GM�p�]�~,�l�?Z7.')�He��R�1����ۑ��lbad#��d�&�~�`=���;�=�S�6I�ܤU�5W�
�4 ������hY����~��/�sc�l��a̢�s�/#4-���13ָ9M�$��*ݍg�T���n���2��3x�/�vh��)��v�����&Y���>�ps�< /D'����+Y�F�ſ�-֣� fj�%����zg#S���X�cOM$��ɼH�,��e��Z�9��uQ�����.�h�!R��`.h6p�"2�:4��ٵ,����lp�B�l����́+<��։	G]t���-�%�f![�uF���31fChn{��Q`FL����Z�벴mp�r5�p9@��h��Y������%�d_�]�ޏ�f֞81u�Ųf�f���Ԭ�9ؐ����ߒ&s�8]f��O�d�9.�2s���s%��v�� i�Y@�L=��1b]q�/���5C�Lx�/�6��Q[Nq��,4ۭ��d�fհ�[?2�[�[>k�i�&<u�ͩ�p�B&z������&Ƹ/�����f�na��ocGe�zk~NL���u�?7���.ƍ����G��^σ3�e��9n7�xܐ�C&Q������q�g�ԉY(݌�31���u����VoM�����&��uw}����Bc��w�Q���m:��p!CB1d�Ժa4���%�˹�j�05{n��n�}^�,��Γ�,�k�;�g;"7{1b�v*�Tܽ�u��lē�PSC�K�N�|����\�����$��������T�W��ua8��$��������p4aJ��̸�r3�
L��;�T͹��ݵ-_-fh�To!��ѳ:j�D���P�{Y��������Yq6շA�
�b�d�S�	��@	B�'L��\y1}�90,�2�r���IΊ�9�_�d 2@�4�Ƈ��� f�\n�>��Y#7I��ԭ`9{f��^�$��\g*3˃���@�y{���B�6r�Bh�l��bs�q��G���2��MF2��z��B���ԭ��ԁqûԿ(u� ����@r�l�jV���i�Z���� �UOo�i��+��p������x�`bT[N�K��d"��ՠy�RG��p�I�F�R<��[Uob��s#���,��j0k=�3`=$,~m�/�e�
�,F2�ds�ŀH��[���YV�$r��e��4��=8+GMx c��̛�L�0%'Ӽwsp�S}�3y��jY�ĨY�� 3�X¿(ur\ܬ��c)�^�9'�'i#f����~�,�8Ç;�躑�.m�ȜeǸ5f>�1p���S�W�	��@	B�'L����0�.`���W�Z�����t`A�f5��#�q� 1S�o��gb��n�v���bf��֚��,�gix����������XWs����c&�~}�@3�br.��M��/3`�l�{|�_L�q�z���T8� ���f�?;b٣����eˢ՝Pf��3I�1��'�#V͙s��S�&G��̹������V:��ul����2]�ʭ�w1��V�͂Cf��R�ŝ\#5pb|��T�:0Q��NLJ�Ø�-\��1�1a3��1IjG���ߜ4��LҲ��gf/��0�m��\8p�D�˲_H��Ä�ꟛ�k�ܓu�p����[8�y����(uhؼe�.I�G�#f���<BҿG&�R5nn������c��%�s�7]x�8!u �
�/O�dY�b�h@_j�.2ky����$g�A�q�ܳS�LA24b�~�Y'^8�v�O��&�!SA&�u�	ſ�uQ�2��-5n�v�W@�.�����S�"�-�+���X)��}s�p�.��fA��u�3`��)���,��as�Ŵ�r�B�2#'��n/����^ǭ*�l��`�lg���������,�mW����uſ#N�=>GF��F�,4�M�ͺ���l�M���m���Y�Մ�r��
3�'�LS)u��fk9�s�&܏RG�BiF�����踏f5���
#p6f� >xJ��jK�̍8pl�hZK1�����$���.˫|��n=ͬ�1�I������j"�eR��ǋ��q�&<�7#���:�S����37o�]�uj��Z���~��*_p6I��<�Yzw�d�[7+/� &���.9�r/9�n4s�,�'������,�U���s���ޕ�jnLwb�\ﺅ���]4I�7�^n�⫣�e~/df�,�ep޸	O�U߼���J����rn��O29I�T�B/������G�[��v4`^	'��DsH���
8+/�/�̯8j��Ǉ!4��uYhn�7�^�#2L���z�yߩ�u�a`ݖ02ɺq_Ί� �:7M��01IDE����8��:�:E���� T�~y�$�W�fEG�+��fl`�ݴ�.�zf�9$1S�b���<�*����Y#7I�E�[�rn��_lb33�tU3P�"s. lȈ�E'< t��	�FNt .�����1�oC8p�1RQ��ʋ�p�R���/J�%8��,���Dz1�x0�P��K�-tr�J�Փu���j�Qs��p�ȹ"g�v�&F�5��+9ꉉXW�?��e�����gsXқ9=u�ι��/M4��f0�,��r07�@���)K���AkYɑæP{e����'A�u`�us&.+9W8i���z�Y��T����mnC1u7I��z�-��j�jS��24�&<�7wW��] �ZrA���j]�Ĩ�䙏�I��Hur�ͅ�FNҺ%�f�$7�F�*�k���C���Y,��,~����[�!C&<�#qL�
�C�p?}�N'D��%�_�0�g���3V��hI.���MK 4��=1�z|�)0JfX�v��%�nE�vf.Q9��b�l�͍�b�U���.̅x��IE�/�NL8����b�#36��^wp��Nh̜ j��IR)޿�uQ�e�M����͹Q���/{6��W��rޱ�n�IE�V��Us���D�23���S�q11N��9R��Z�����5Xg05��u����I��uu�@.A6h��}U7�q4�/��0թY�巬r8j��G��R�*m�n+�&�~Ȝe����4�׃���1s�/�d��.,�k,�}ݩ6���m�$�[�����u_Wg%�"��olN����9kj�rܴ��#�LJ�I~�]�}2@ם����#'ة�~\��P����l~y�I�w���=��:3r���S�G1�]pnV��T�/6�h͗���]�M����YW5��q=ƺ�h�𗀛0aky�ܶk|.��a�c���͸�Wח�u_������y�ֲ�̬ə΢Q�������M��������M����|x�����ˊ0oI�w#�"9�^��u%����5��FY�Zb�P��U^�g�21��zMn�C./2�;�94F�D��2orY,
1밮bj�)|b-fbл��k�@v�b\��h1�{R�C�I�p����5�+w6���Hu[ދeq�c�Twf^��3	g �3f�,����v��sƸ}Z^�-fu䨉X>G*S�	��@	B�'L����>�p3���Y�,LˆMm�sΠ�8�x�� 1S�9�,L�CB�t�.\��{��pie��Ꟃjؐ	���e���z�HK�E�/Z]�Ԅ�a��bw3v��g�cg]�$�x��YI4r��+Vn�{p��b&�`��g�r@]�	�q_ż�LϙM����^Me��s���^3Ix�T�5j�m-z8h�TD�(G
�S9�͡���-7]gf-�u\�ۗL�Gf����6p[�$F��8���U#'b]I�l͠!�"�b��D���d��Y��w&.�l�Z.����;8�qs�_'1)�"�m����4�)�^wܺY�n�-0�n��\�bа*'�_���n����LN�u�t1�W��R�f�	�Ʒ�\�Ka��)eG�:���LLr3b_j��j���]{��O&LUb�M����R7R���܋[��Ĩbf����p�45%7f%Nx3rb�<<����v����=�6�$�n���:v�t�s��+GN	�,��[���MĲ�_�b�p*�EO�lѬ�q!��u��[b�����]���cN5Ν#s�3�&<ul��}8�N�����\ڥr���z6�o�HY53����R�F�5;�R���!��{���s�:��Mɉ��(u���=���:���F�ˀL�-�%6L?���Y�1�(�7�ʲ_hV}�.Y9#��^vk7`����#w�%~��S�B�C��и6p�>E([ً�+��M���7��ZA@��l1�!���1c(��ty�9<��X�}s���u^�nȐ	S�(�t3p�T��I�r�͜���ꋩ�Gss^w��I�?����רA���
XJϹ�E'�A��a�sxZ��e�&b]�25j��2rVD��0���n��x���Ľ��x�O�=�����dC�(uf�l���61d_>n�@�&ח����uV�%�8zlf�G��c&b]���h�ޱ-,�p�̙��ܚM��"N�@mJ*H�<a����� �<��������lͰ�MrV|4�~eȸY��rB��GC6���{)�9�f�I�Z�ۻ"���
>�떭��ϕƕ5�58��I���܀%��,{2U2��T���"�qV��J�74f
w���Gf�@¯W-��S���V �eq�� ��ͬ��nj�e�|���a(�OĺQ�e+g���vĺm�A��X71���/��]�fѲ����L���-�5=��`�D���-�u�s�1��9�K��)zH@�������ٞ4~�oګ,1bj����x,11,^e2ˎ���T��W�*f#b6��[�ι��r��Kl����.Uүg^Ж�R���$p��`N�j/��7`���Z��+`e/�͍���x Y��%&b]ʩ�/�S����+���?�ߩ�3��&-�$�٘y�E�ƌ�b�&Ԭ��̆�l=�%0K��%܎RFfI,'6WQ3��������i�[�CՁLRH7j0�b�T!���#�X9"��@5�
�𵪴��sM�Ӡ9FH�bu�,O4l��z��*.�#'Y���X��BS���Gh�r�"����J���qBj;P�PA��	�, +t�� �e`�Px��ܘ5@��6-ޅy��`j����f�r���=:'�0$p��j�d�^v�]��%�u���+u�G
�Sw��3�]vN��Wd�t
~/[��e��,�b�on�\��BLʒW���.��qI��T�}y�M��-�p�]�2r6��j�T7�|]�,Pۥ��X�*rnɫ�	����]��LL�uXRdn�t�b?�T�Ii�����R�p*�n����f�ϸW�����6U���W��M�hN.1�%6�?5g�2X�3���c݀�9Kh=�l�_Y8�uE�:��-��_-5��%W�9���aE�[�z�-��NLҷu'��l3��������r����,!9�jeW׌���̃�:��48�Y����x[)�̑�,���u�4C���(���u9������bV��b'��8t��2Y4p&^M����xY	2jb����㮘j��C�9��u�q?�n֕XJ�Wl�I�l���*���1�L�ĸ�f9�9ȍ���|M�As�K�k��X�`ևLĺ���]�n�M�1aJ.fX��Co���f��/E��n�����Y!b�$}�R��fA�f��C�ü����-�����Y�ۤ2q��Y��;��A�.��	6��TM��/70h��k�Km��c&�~����0p�o�[�7��$4�c5��2p�d��p5⬓s�^�G���u�uK}Y�Ȓ8Ô�8�0�,pס���9�����Dx���i�� ùud�p��� i)���W`Zxg�_��wEc�6�����D�K�7s���S��0�_?4�5b�ur�������M�S�	��@	B�'L��\�>�p9n�r�͂#f�)ݴ��9~Va���g��v�d�� fb7��;�Vk�.;1I���I~�bs��J��!β?�$�����6wIL�ԝef��Y��HM�UQ��VE.8!(׺�a0j6����j�ĺ�غ��L�ԭЃ��͓9R�ZG�/�NLX�6���b0뼌��_���+�a�0!ȷ��!s��g����}�AC�6�Rw��T��0I�м��/V8Ӯ��f��	}4$�u	�>��ڋSd�V}�_�[�q��c��܈���,�viVJ�2��&9���gi���b��VТY��6���k1/��11�_���>H���D�4�H�F�3��؄���i��qc�mps�Y^rק�0���`�$��B(�\5n"֥,'s�m`m����W���[
+����f6�p�Yt�M�0Ս�l�+�����E�?
��Yce�A�;�{�pX۷^f���Q�&���-�g=�ުp�]	6Wd[7ͷ�E�4�, �F&	����7�\��;.�ϛ����/2�z�٘i�V��h3`�,0I��7��Y0�#���+`%�?���#&L��ʬۦ�ؐ��/\?��l$��k�<]13hj��{@~�&b�/O0h��:Z�Zk~<,��7C&���t�]ݕ)r���Җ��$�Lfu����2�H�t���wY���ۚ����`�j�������&���{��Y)6b"�e���I��L��/m6��i�pW4�y�������$Ah� ���*��YW9f��E);`�3�*��I��R����,��t}���R%���n�̀�o�f71�=��.j8h䨉X�U�<2Є'=��C�F�!���
�p.+�C-�CY�.
�9�ޅeQ�IZ���f�+��	�Ռ�[6`ں���T��5����{�����_Z1����Ⱦ����B�kB߻Ux�[Sf������i��R�X�s��� MxR/u5�ew�k/��p=�����L��:4rn��#sx�Ig�d�Š1C&�:�8!�(A� ��I5Gs`�\pk��<��cn��6�iz�9���bb�p�҂���BV5��(���&	�7h����l���U=�Vf�O֡y�����\��.��*I4`Vn��nv��<�9O�$���.�c��%�3#�J/��KS����fu�T�N4ۮß��`6v"���&�8i�܊SCM�NtȸLl�+���-=7�n���iq!E��g�$���4"�f��NQ�<wkI����;ٟ�4� �B7w@^�1�s�_�p�,0ח� t[�Tv~oww�%�&J�]~���z�ƨ�N͙��-s8I$�!�A5��i��sh�`�l]��aQ��"3(k� �Q�&��X̆/��	W����ik�L�[��8�&�e6n�p�^NO1Wi�t1ɉ�����6�b��T���ohbd^����/p�r�H�*�9��P�@�Ý~տ�2s"���!��hQs�Oj*�DҺ�^�f�"�e�9i��������&�9�#Ma��9��!�&�^�:7l�x�sAL�F�[��D�x��j���q�fI-1�_�d&R����[��,x���^�5��;F�C�*�Y�mk���u87b8���Y�5�����11db�� �m��qS�gV+���a����͕*1���03<+b�����z�!C�p�;Mݜ@]�樼�g61$[�����a}�D�K��8����",z������N�3guV�Rؔ�$��%v>l|Q�)�=�1|j?@X�[VjN�զ�X;T�鉻��T�Ow2ǚ��������8̨��Zr�<۝�A��4K��T��Qs�Ԡ�GC���j.{1`��]�e6F�ȿ�/�+l�`M�W���L�E��0Ԙi�b܏R����������Q�[��wcbN01t[8�V3��ÉV���(��qs��d0��ڍ9�%�*�A��w]O���x/M0j� �a7qh�@�U>�(�����"Pہ�
�/O�dA�f���eqL�Y�N���6hj���LE����|�9���[ĕsA�h*����Ml�é��]Y5�}w�`��}�/�ўL�k��9ɜ�b�$[�����*d
w�}e��Yפl����`1d"�e�3��z��,�0�_���y��h*��,�G_nN�d�&����֑9b�B��z�����{�|�)��huO.g�\y3���ݹ�\�S!�1qg�9f�d���������f�|2Y��|eO�ͫQ�L�nw��7l*�ޓ�ֲqù{.�<���'#f�O�8b&�v���juיY�#q���n���e�8�$��T��d���^}81�˹��و���Z��+���}Ըqs��L����C���M��kS+��n�D,K�ڍ�C�5f#'L�O�u_`����r�ơ��c9ב�13���c�L�s#�)�����upN�%�fy�>G11��L���	� �c�
��9)"[�� �����u���J�V��l�9�V�T"C�����p�l�Ĥ__3��K��X���b�/�k#����z��3�rz5n��+�FLԺ����9�rd�T��sῢ�-Luj�ȑs����$��Tgf9/�C4�8��t��zh<��:0�p�ԨY61֩�,8�g%�zG7l��e'F�����zp
�Ѡ916� �S�z\��|�^�+�ޯ��?�[�f��-&S���>1Wg�IY?�Ss��Y�-�_N+�f�@&�~��ݥ'f�|,g�#��-jΠ�#���^x�|Y�`��UZl�֋�LK���������<ǦѼ�M �YV��aЀ�.���l�mk�14�I�i4'��~=j��3�{C�L'D��%�_�0���}����<��Nͤ�Mmb����܄U�s�b�j}�z7ʆ4���U3�2�ME�R�>���[�+�b����Gws�H9�F�&�\�.^�f��#g�eb�M���&�p�꺭ê�� �fY��8��$��9ݏ���)0��>��<Ƨ����#f��Q�,c3p�<���u:�=��'��&n�&���4T��Z����f�%q��$�@��l�D�g�x��V��q8]'7UD6`^r=��I2�<����j���e	��۹\����)\t��X4)<��"�%4+N9d�lv#���'�G�3#F��/�����M`"�-�g�毝���+��u[��ZwF.5�z6�d�B�.KeS`n+�H|*�����A��p��z��� ��tX�.Tƽ[15���li��d܄�N�z��RID�[?4WbE�K��"�Y7�����cr��y�5N�p��.0l�(]>+�2x�$x�=�6bq�l��R_
����Z�gU	k;�J�f�bȈQg��뫶��ϟ$\���5�Q���"��y5�V��8��ܹ���k�&��@��Ŝ$ss�k݉�,��g�16����%GNC�Yt�Ww(�&YwX�#�<���X��~ٜ,\_4n��������a�t[jFX�<�$	~����"s����y���f哪E)��!�]���u[�9�.�N�칲j��qs�Vz��wn���j����Q�h*��6��Pw@J�<B����?�W�P������۵��7���,��.���#��9!��ɵn��%Ǧ�(�Dk&�n�5O�o:��oQ��<��Mʁ� ��́�����祘+�o6�`���w�.��Ы!CF�%!'\�p�,=���>�RV��B1�2sH���_�hVg��i1����'�#���7�N�������FM�j������.��C����A�,'�6�Ӎ������]>b��Y�b�Sw�V΂���t]�-J�!{3���L����L�M%����m�r2jN1rd9Q�,_P�,�eu�	K�H�*k��q���:E���� T�~y�$���~�Ჺ�O�6G2b*[��bm�����f����ɂ�f�C���ȩp���Yg0�IM��s�>�#8!RwY��hS�8Y�0]��YܸASA���xeH7�9r6��ܯ��Y߅o�m�M�lA8��ܺ.\p"�e�.�$�n�Q����e];6��r��-1b�$q��`�%��n�Dx_��q��T�9��s��Ǥ�����"�4L�o~ch�"��B#'�uٿ{�����K&L��4�!��c��s<�3�0�M�p�#GN����ߴ��F�d5����x��m�p\�e�f	�	O�����؉#�+��꘩$9b�ꗬ�! �x��alOL�S3��������r>�����u9���9_Oǅ�L��?��T#fmȰ�B!s�6	������T��"�E������u��Fفa��,\d6�� 6d���Cf�%���РfQmY8�<r�RҚ�1��p��Ű)��|���b�$ӟoϸ�p
�#e]7�|W�_p�ÑH�.�R��0�wsX?�5r
���9nĄ��̉�|�\q91�E���_5bV�8既��e�8!�(A� ��I3ס0\N34fn횪Y+1d���г12l�l|o�����K�l07l*�����b0�ln��+g5Ŭ���[ ���'�^'��Z��:�S!a�,n�LeK������Ƞ���Y��g�3&��w5Ĭκo@Lĺ�9r�s�a'<�O���sæZ�4��-FL[���,!0�B͂�FNx�������f*a�,�-�,��-i�&���3q{8rȄ��M��r�_72r�d�>KqY_76�I�18�mA'�6\�l�mY�uF�:4`N���r�$��R�bn��	f6a��(u+�r	ރ&	9���ս9���m,�l��bȔ28g�kVzc��jN�U��Z�Dש��5z�81���<*�A��Rz-k8�k�Σ0%_���9���)����8����g�絋�/B]ta���p1�a�w��e�f�,�d����(ef����c��L����C���¡�����ly�@8��-7T!�z� 9+�P�Q�L8\�cn����j��+O�FLx8vA�YH�Ռ6+<�����_�n�]�h�nĄ�n!9�ݠA�4���_�/�%�f�ŸaC&S�	��@	B�'L��� �e�Ac��������X��ս�r6��l����`��9�f��iَ��|1��^6�51\N��uS�x�Tw�ߐ���QSХ�r��ꬕ�d��[�]8��	�p���ʮ/3a��>-��=6�T����g]�q�ϼe�2r���v}��A0a��h��9X�i;11u�29�����M��9]�)�0����ӟJkS���H�r�Z�G�����%*�2zA^��tŘI��*�͋b�9���"ud�'�bf�`�I�-{5`�#��L�x<[�%�)5)���ί�eT��M�U_V�5A��d��X�]5W���ߺ�YE8K'Ʒec�y���,C5ɺgu����u��\�f󇗤_]�n6��W��r���N�Y�}�n�Vy�Xw3p��780�x>���ݷ���Q���@���]�c&\��P�aj��PfJ�	��ً� ���p�ð�a����U#3,JYt�-7���14ab�*�<3�сFMx���.��_w1j��݂�zbƖ*���ɍ�lfl��\�M,)7+7P*u�Z�e�`4a�[�d�y'�6	�_p��BOƌ���5�eM����d�9���y9pԐ�:6��c�L� Q�?���Yp�E�Ҫ�T;�.�9���	d&�e5hV�"��0�T��Aˏ�nw7�]1�����{$�F�����A�.�j�l`}L9Ũ讁Y��č6pЄ��K�.��c���"_g���a��Aom/���}�E�vl�r-�6n����Va�j:bVp�fN��V�M�sf�7<5���E;��r�S����x�#����|ln��$��Pv ��r�|�I}�#���AS�uY�7�rf�$�Ѐ1����u�X��ZNn�Y��:�Ô��\6rԐ9kk�%u�5�f�*Y���k�/녱�?�ӯ����1,U�f�v���u]:�΍1`Ш��zB7�w6r��k9�gQ��a�ɿL�˴�t/���6�[�Ӧ����4{b�lL��Y�,����'��,�����32n�49�.��*��]�5]��<��j�!��������3�9~�$E�TwH�	'�2��p;J�mɰ���n�M-g�R]d^,��o�S�����:b��ٓ�Hf��z��!���[O6�$����!i�����ҳ.���"3�ze���	1��:4�|��sɚu��X�+�f��c�q=�Zw5l��)��v�����&Y@�c�� �e����ct��AS���= �F���]�ڛ)���w�as�W���Z�r+7	�����Evc�M���o��#�%�r���p�Su��7׶r�E��yLݫ���Z��.��vpԐI�eC�}5jN�L�3�/�'����&�A��q�.���:BO��~��d�<�RZ�G}��z��`���
?���n�lj��sEO�d�k�7d4�M#�@���Q�������|c���qM�u��{}��1�.����Z�d�'�z��(����u���d���hΙ7��d����ׅ��f�ovq}���+{����f����?9�d-�~��(B���O�C4�Ol�����Acq��빙���;ƪ���u1�19M*1K`I/n�}K
��;&��.��m� 6�=\�/���B~~T��,I5;F�_v�r����+B٦����51>-��'���UZ@��tX�+G����{4�&b]�mٜ�o\Q�R�`��a��AS�֍͝�������M]b7�4�u�9���(���{<�8GC�������{O2��=+�Np2`<��Fݘ) ��"Pہ�
�/O�dY�u��%fj�`5�~꠩MlN3���/�;��5�"�3AW��"�2Ws=�7�T��Z
n�[��>܄H�Y�eK}��I�z�҂����U��sڲqCf*�d�^�fs�"�&�/�n���p�:4�Z�a��E�&b]��̪.�cd�0�.䏵V/��ˢ`#F���US��,���M��߬��Ϊ-�ʪ{v��fb��3�X]`�����Jf�v��ů&<�_�e��!{b~٭��as�©�vspC�Q9g
W���:�Yr�,����l~ګ���$�.�%@��ƶ�"u+|�ts	γM��n�lN:6qB[=1CB4�d�?3^sL���|��Sy�p��+3l�8���=Ȭ<��u9�9�5h,1�I/�:m|�G�,42��&ˉ��(u'�E�p�Y�I���E���{0 #�-ߣ�-k7�x�۬�DE)3����Y�+��L��o]�'3�Sn�͵;��XvE7�ͭ��֭76rVn�&�&�~�Ԍ�l�B��Bc���F��q����h_�9�&L��,��,�@u��rn���cWL��У}y� 1rb��P��b��!#��X\fܨ1�)��v�����&Y@�H=��2Xg6l�'2pAO7�Y��Fe�����w�E�5�,��9�r��>����G�ں_�!�A�L�*,延F�:���ٚ�/B1l��B���O�v�̨Y����2]�X6y^}[�d�-8�)7g���b�9p�'�6gF��+�� j]q}��sܮ�mF��� ��n�,��h㺜3~Z�[�,;����v�U����ԢX�[xʖݙ���2k��D�[��=J�BN��뷘�o��ۚ���G��8��7ɳ����������j�9?7rUr��ϵ���B�&Q��nrٟ`�TهRk �� ���ହ���Ԫ-��2a�b�$�N~0ߺ�9j�s_̼:�ʫ��n�'c�-;��A��ȿdj��W��Y$�E9Uh�eaYǕ��Lφ�@�J���K����n�b�v�Yׅ�}f"�e�Y�l��v#&L���&p��jF�dj9�����U��6�\91��Q�����Ą'�z�y�몆��d��7���rtE�L��f�N�٨�X�}[~d�bf`Ȅ'�*�o�"�x�o�90��EfE���� T�~y�$6�́�les[���}6��z�A�Z��Ts���t��:.�84m�8���*i{�:2?Ϣc�M\,����c�Mx c��2��͸� #�(��_+'<�����@&�����m�dY��U]��sp�sN��������̷�c3@u�>�4���_��/�c%��!r5�}�����rts�X���8�����lC������v�[�b؄'���f��l�2U������d]֟g� �ʛ�fH[�;-�P�S��f���OR=J���Y*�t�'��|��U���t��k`栵�l��t��/���Hu&�"s����Z�:[�Ys3a*�f}��E��\K��n=�\֛YjrĘI�?\-,K��ӈ:6�D�7+&�?9�Ofe�qߌ��uYh���.p�>
�ɴJK�(tR�	��@	B�'L���iF� ��.��B�`�.����ڴ���Ɍ�d�,@��������5�\��A�3�2��"g�yؾp�Rud��U]g5+�&Z��R�\Wu�+s���+�ͺ-��:7'*��a3�^�XH��<\�pb�?�s}*����:�y�]1)�E�{�U^����E�sX77f�V������1�-0]�$�\��lJ��Хr��ȉ��,�7KLC���up�9���P�U7`��1���ӲU�J3d�n��9�@������T&*]"ԉI���BfA\�h*��r6g�'8d�$��n`=���(i�4�캺��Tw�e��D,���(?'�,��3g87��[��x�X��r6{�^w71|�P��΁euF�1��g|��'c�mz�/��;����1��u��ج65х`C@�����k�����1�*h�bB�,:����.�1fBѠG�f��yR:\_�����p�E�scf����h��Q*f-98j��H�ӈ�28��,�d� F� 0j�tݭu���pi�1�����[�_d����0vҨQ��I�v��s�@#&b]��y%n�Ñ�+{$��:�y�C�&��[6�y!��i��/2��A�Mxʖ��i���&	UQ�F&7�;�&	0K���Z���x=u����a�((Z����J��A�� �_�ϚT�f����z���fΧ�U��WJM�p�k|��X�I�f�p��z��Lx�/[0��uܲ�����,FLR�5Z�C؂�f�5U����*8�X�l�fN�]9�c�ðYHnG��'��c�0�N�z�Ya���Թ9ߗ��f�m��9��I�����}�n���'[�G�#���f���2��2��JG�,,����%u��j�O�
��M��*E�;A�\ �7r�G�[��[�g�B���`7n���]�r��<ʥ'#&���v9bVT���uYH+wРy_����]T�N'K�� �وA�D���g#�q?k��!�'9[%�nK4��.hLq]'D��%�_�0��*���}�ڪ�1p��~vӣ�&2۟�˙35��q��<�Z�E�&�x �L�_Q�ȘY��/]�01���݆���{x cIoz�99*.���.r����,2v�u�.�1�������c� �hu�����E�A%�_�����7�I��6�vۘ�u�+���[��+HͰ������жa� ƨu :6)g��D�+�g ���`4�I��s��$s8DS]�kpĜ��d]V�[�M���X�!e��]��~�Ā�S���ky�b���`�ܓ�>��� 0`�:�SMץfѺY�5���䚾�2EX�u���w�հq��f2�DK�:6�fQ��������3a*3���7{�'}�P�bn�7�',�\^n�T�٬���#&���:�߂ �Lĺ,,6�gA��f̠	S��&��,�Q��)��v�����&Y@Vm���:�W��R�䖔���4��jc��Ɨ� 13��pq����ޘ�F�F��l�I���M���3��M׭�i�y5�21u���~`^�u�F�m��	��z0g��Y拿�VT��1�E�&E���`%߻�#b]�oU7}xx�6�I�fA��C&���,�u���S���yN��9I�#՝��o�fR }6�3s��t�}qs(X۵��ur6�<Ϋ�L׭(5�Ȏ��I�V 9�:-�5�����=@�&Ʒ��^�N͚�/_�fb,B�Y��gc�֭�h����Ki��'c�#s��͡�_��*ʖ�Z�Q��/B�e�s����$��\�2/Y��Բ%��b�-9�,i��E�ɇY��]N׭������R-�����X�I�f`B̶W8j]N��� sw�&���v��l��r�T�/�Ӓ���ܠY�y��.�nS�u���.[���;p,U11�ǃ�r|��('�n��yǩ���b�f�&���U�`��8�����U3�%�u*��m�<���uٿ������%c&L��v�ą������Hr�JG����m4� '�_�:2W����LLˁG���j��������ag���4�Vĺ��y~�v;7�J�7v-ĸY�5�F�i��H�G�f���UC����`}`ԈIB�9���{f* ݨ���B0q�K��+kMĺ�c�
+vN������w��������3�-�$G�[�͝~��NE([:+��{HdΪ[�:dȴ��m�������c��\h��u&NĺTv2j�\���a�&L�W��v��Mu�,����qBj;P�PA��	�, O�.��ټ�b�Y;1'/���f��:��qV1S|.�%���SRm��\�I ]��p�9x��!R'f2C6n��Dݲ_��a0O�FM�ԙ�l�$�5d��E�,RYy���<�}Ё�F̸k&<ڞH�Z6�Rwfn����Z�Im��W'&,u`ܠq�����ᯋ̟(���?�5��n���b���qt{�j����]�22n䬃0㋛d��fP�FL�������L�uK���݀���ʱ��m����|�d�3]����_d�%z?�Ո	Sr3��)o�3�8hn�(�&��(u��h�c&�[��Ȍz(6�V[Lxh�j9��{��Ix�V��#��M��nn6��/��[�`��D8�:9�����D�KY�ɕ9��,7�Iof�b��!h�b�T��\8ws���n�~1�u��T)J]dy# 3�P�!e`������x�{~/�	K&���fx�f7d�T����3[텳�7gAts?rߗ����!�a�ߓ���>dn#g��+nV�Am��?�$r���{��Y8+�D���ͼ�<\8fԄ)��ܘ��Y1M�~^m���&�}2r�u�脭u��I~�c�/��ؘ�f�hj�s5��6��`���9{���E��j�IR���Ȧ�Yb��bοShS+M�L�+�K���T�������L����~Yn'FMĺ������Z�)�z�$'�
�;H���ȐI��oSwYպg8��R�	Oݪ�,���M��HuKs�w��մr	�/�%�a8��ԭ��.����`�^�d�c4r"֥t;K���Q'<��z.�C��CL�����f�x�d]0:o��S����u�ꖵ8�y��oH��:�ݦ�[�l6=�]�8օ���Mc�YlN,4�3�O�5\�]9���Zfd��g4IΝd��ж�䨉X��qa���	Sz6'�kĀ������`��80c�c�-+u�\��]pb��9�7kg���)��v�����&Y@Լ�0\.��L�z4�A�8;M�+�fq/8�3����ͣo�k�k`n�;�,19I�f3T�Cf�UE�뺱�&�]�N��v��lh~���=)�q������=��~�^.���+[�x� S�z�9r�\�%�~&8��x�S}[�5]��/�.��&�~���Za��c��/g��&�ĆˁJ�S��NxҿN�%�����,��9��,h�H��H\��s��!S��́Q��&��m`�ޗ��l�mӻbސH�����)n�`�SpR�"�ݭuRsf�QC&�[��e榱Y��'F�(u�ǫ��"w��s�̴j��$g�vr��`��cLS�l��¶8�Ĺ~���kw��	S���1u�Բ��r>7�I��Dέ��S�s]�ϡH��8�C�v��a���j�f��� C��ʮ�B@��'s���e)'�ʧ�0b�m���o#r����$s��1��Է��Y	�Lj���C�zf@�P�S�Ľ'��l|�\'5n�Gof�GfĤjE�ss�T�ɳ	NHF�;�U٬�9������9\�i��y7f�tB��ܲu�s8�h=�=p"�Ĩ�CfV��_���Z�e����9�W�����!��`Μ����fn�LOS�e���hbX�(�XWj�n�Ժ�К.�m��@K����1pe�!ƿp��l4n�nkf��31�Q��5\75.��8�ݸ13 ��/��Y�j�2�ݻ���P�&�\̙zt.��Y�bsf�Nk��aQ熮�b8�ԤXc�<����Tk�Z߄c�\�1x�o�-��:0�}n���AȒfg�X�CcM���/{3�v�c�g� �ąL�ʺHdb�ɧ���PM~�:Ԭ��� ��upƇ�n�ĸ���}[e5+"�ML���ߺ]�u�h�u`Ԭۊ\�� b]�z���gH����jN��R�
��于���&<�sPxғN�tF�ש�.+�未n+��v�����&Y@�n}��٧����ǧ����t�c��q7Cq fjh8;��-�jв���fSK�G�悇��\�v�W�L���]��|5�Y��|��k4v�A뾩��GO�;�D�Z�9����@��s[܈�X���9r~��<�\��.������a0����f�ߢ�̑����m~΁uT��]�smM6�I2nbܿr+�L���ʢe{�l�y�$ɻ ��=�հ� "f]�h�R7�ֲ~8jN�hu�c��B��6�I�ʛ���f��G�
q#�Q��t�-����O��\�Ű�KUM��p�!�{�_ˮ���/��:��T[��Gf��f�\ ٜ��g'�p����"֥,>����z}Є)���YX���s��wp����,��������j�*1�~�9×���C�(u/Xl��J�IBn��s�l�M[\�D���qt�����e܌fb܇�f�.�C���.4'�2��f�'=���NG�vUxg�̀9���o��f�<Tw�5�ji���$��BYW97����*J��������8]�����r�U����5����eၓ�_���������@��pN��\��E#����n��\��ԑ9�ݜ�K�$v"�~6{d�Yzn����M�����
i�hܐ��M�ᇖ����&b]6~X&���)}Z�47�L�E���� T�~y�$��f�0\��h3jV��Y{1�6��jc'�Ɨ�6jֲ_w1l�<�"S��̗��ɬ�8I�,��X�؀9\V8	��a�,#5��l�uw���x�S�r�_�5M�iћ9����H+��t��,��#�r�����[�f"�e����f��0��Db�̸S|@"��F۪R�F�����z��2�1��v��v�)^�e%*��7y��k+GMx\Gs�Y��u���jY��B�%+�r��)���f��%aS�f��,�[���S���lj�,�j��E�[o3�t]o#�d�����9��&4�Μ%��%�fc���%��q�a�֙��r�(�B"2j�lլ�$'&�*L�m6T�s��B=��I��g��]�Jĺ�N/3n��'L�r�������8GBa#����(H91�E��,,5f��Y�l��+a�_v�Zv�2�*4a�CfA:<,���}7G�CCUg9�9�/5�X��W~�
$Xѐ�����d��Ӑ|��	�p�n�A�ii&<�Y�ݠ9�Wl�W�Cz6�p�ש �Z,�v3b�e���u��9~c��P��l�\+9r�<	��R�	��@	B�'L���y�>�p��8?���Y-4hj�j�����t/<kYC��k*�BY����0ɬ���"uk)�Yǅ�^!Rw�=5G#7l�u�v�uf�������@H&I�5��������k�뚊I��k4bn�neM�����'��G���G�1`6,gLG9����Z��$��{CW��~d���ܬ�����Y����Y�I��,���ٰ�
ap��8����Ve�6�<���5�I/�88 �Q3�Ү�o�-u#N��Ь�I�Q3�WM¿(u���^#��]̈́F�c.8�����K��ܜ$��a�!�$͈YB�4dԀ�J��u]��K�_]6r6��`����7fF2��jĜdǢ6Q�r�`��a�,�	S��97���BZaK�o!���܋���c|�PYHfn͙?:�	��n���3�4a�CfދC!��3�빁Zw>/H�@6��mn=N��N�D5[��`�,�7$�/�պ���B��BZ��]�m�A#&<��R^���ZL��0�G��60���Z�'�
VcFM����P��"�E���X�FĈ!�S�8!�(A� ��IֺK}������f1n|4�i�V�8���f�)@f�����VN�d�2:oȬ�y�pk�� #��j�Y�a�3�Rak��e}�̀�2���*5۬���.���#�m7-L���u}�G�|��I+'&���q�ֳSNX�s����,{0��(��y�S�L�-���vrt8aI�*k�>�p�tx|bs���d�<�D72Ą�pq��H���Tnj��[m4	��E�{]/h1�q4r�,��3Z9��y����I֝m1gK6`*ѯ�@s��x_��%�B�MW-�����搙�ؘ9|��&'V�fKme7����F([��ֱ�N+��d1�ͷ�>-�e�,��&����i���&Vf�r���ݺ/��̝IցYAϪ����D�cp`�庉������0.J]d\��pῒ�aX���b3q_V�Sxun�����01L�s#�j�Y�.'7�a`���\~d���\�01�%��� ƍ��0t����=ԋQ����b�d6�fp�\���a����	�:1�r�ll�/�5<u�1rή��$�^��ZͰэ9S�rV�Hw�$�έ�]0.�g�N��v��4ɚ(��rScC�Yc���y1_���+hI��/#u��Sdف�67Ϙ%�Gg|�	1�	�Gq9RY�-�d��^~Al��
�K`��n�	W�Ɨ��>��i�_֭�W8�$<�Y��s7�l��\by1�#�M�,[??�E	G�UAia��.{hV#I�����it�t����f���4?[ߡf��ܻ�����.<uf�}O�$�D*���-T��d�:g�-o�̼β_�'O"����p/8/���.���Rsؑ�&L���m��)�}5n��F��ꛉ�;b���e����v�m�11�~�!s<pQ�p g�Nܘ�cpuW���ԫ�^h��Bz�Űΐ��&W�L��f=g��9K6�Z�G��Z�NK��`�z�6-�]2b�֥�!��mW-<��c�d2��g�Q�I�b��,<��ڬZ1��Ű��LR(��Nn5f���@G���~!��B�8p68P�]EĪޚ����7���j��#�6�����Z��1ЁfY/ϵ]N`j�����8�]�M��]����ӧ�_��8�J4��v�f�}����3*�x0Gԅ�N�:E���� T�~y�$��.`�<������fd�AS������q�pn��fJp3g�<@�1S���)2����k��H�R5�&T��Q[@��$�����8��$8a�3f�i����T��u����bҟ�j0�TM�[o9��a�M�o��ɸ�ꭽ���W�u_:db�����/>1n"�e�6���Z��Q��d��0_�o1l��vaI�G��_�K���&�_w߷Z�}��w��-.Iø5�)f��ܙ�N'4�rrV����f�����pb�?
�+{�#֥�[�'���;|�%���ڲ�p�܉�[�pΡ9{c�|�������ֱ13j���L֩Y39WO��쾛�^�CԂ�Tﰲ�j~r�����L��Ρu��9L7��"�愈)[�����d��i	/ӛ��lh��$b�f������2]��@NҲ���9�����u�nn6Ɇ���|W��ti�9��ћ���>�c�_��d�����_��e��o�9=Kh�<��S����za����m�Ñ�&b]
8�4b�Q�2K��=��>�AS��-�����̉��B��RO���\���y8'��L5|-l܈���,�+�.��e�Ď�cTN!�"N�@mJ*H�<a���+�0\�׀�
��ar!�����;�7~�ŨY����ňW���͊as��xR�EI��Fs�x��]��>.���l�g��Ps���S'�ż�"랐�P���USl�d;�6�f��pqx_.ƶO�.��nw���M��_=4r�Ϡ���f�|��n��Zv[��-F5�0�Uds�l܍4�U��f���/s������	��[��q]ȰAղ��t��s5G~����s���v��z/���rR8�X�f���97��E�[o3G���[2ɲ�^�p����	������%W�x	�9M6�&FXjĀa���B"2j6{��:�I����K� G�Zw^&/	�dz8��{}���R:m��^�n؀��C���+ۙӫ�Ԭ����6B�ɾ��9m䤾E��(���%bf�V뚅����W�N�±6�&Luh�_b�C��8W9k(ƍ3������8�6&f=�9�d�Y���.c8r��՜0���:E��U\��Mݒ<��THC��g)��(sh��9EŨ1�&Lu���;N�M��"�]�mଡ7bN��e�8!�(A� ��I3'p`N[0pج����r�c�����^R��`Z3MF�D��YqD�927q��Y3��M
�SfҞn�@�m�qԬ�گ�d���}�����
���}P��{]d����@w C���;��n�O��:7{�Y�ʢ�*-���D��; n`��9��D�+�m�,�u�fj~�Ϥ#y!_����so'��N���D5'��bM�[���<i�:1+�ͽ]dܴ�`�בYN������c�_���p�p6�/t3��c�����<,�:Z]��if�S�쏝�_(��r�.4h:�2Zl��&Ȥ0�t[�V���Ŷ]w�]�5��܈�o9o��*-����6��u���-;-݈1��_��;�Z��Vi��96��=Y �@��d��[����L-[�����821���V�X^���ҩ9Wv�qBSsޟ��*&j]��[&W�Ʉ'�qp��64GM��2�>It���f�K�΋YZ�17���МY�ZKMxR�9`/直l�$Ѻ4N�uGs��)��f�_�����w��ܰ5n"�eu6��r���`���C�������i1�_dU�	��@	B�'L��}� s�և!3`����q�$g�9��?t.2@�����y���`��s�=�en�vG�[����y����5X�k�Ɉ���4���d3��c[�q�ȏ��$_��y�m�~�)H�sI�,�{��G]~d���<6I��Rw����b�[�����s"u�g�� ��N�ݣS� ��c8.G��Z<�H�joY�f�\57l"����r�ͰYY0n~�b��3�Bn1�
^�5Z�dYV_�!�A{P���
+�<Ŝ�f
uW������V��=���W0�$#�!&6၃SuC�RMT�TusIj三
~���}!w3���ur���jU�Ĩ��fPn&�[�:9n��c'�� ���C�!�X�hf�'�b�5\Ω��W�JG���Bs��/��0���!9K����rSW�	��@	B�'L����0�.`n��\rr� �I����
�1SC� 1�ef�Y�ux]X��Q��Iꬎ���:nĄ�n�nb��B�&b]uģ��n��Ѩ���X�tb�u���e"L�k����p�$�n��ew9�Z68��C3�!LeK�е�2QC�L�,Z�9{&\<8pИI��&j��uY\�K}&�ˉ�;0��Bz��s1o�Բds�Ьt��'Ӻ���+Y����+`Y�9�B{�7�v5�ة�f��j�$��±Hu`��-B��Կ�,Օ^ln
����Y�󂍘����x¶�1ֱ��Sw՗k��.�x��b9Q�g��,ۓs��	N�s��@yh�&)����긄�@,̀�����G�C�t�l�}]	�G�#s��j�<B��X�(Ό^�7d"ʟ��ܢ��q]x�8!�(A� ��I�ӱ��5>���Zޤ�6�Y0ѠJ�i7��LA6�u�39h�	��&�s��dB�.:�����5�i`J�M�as���m�T�/�幚oD�&�B��S�����}-�6.�;dfc�Le����ɲ�۫IP|e��ſ�o,uKx��Q#�T&��[���qsyؘi>L��]�5����uj�6GҒ���yb9�49I��Y�՛�]65��D����_�1u�텽�d�T�on���r�����1s�����̍�EUc\W�����PSj���<asֳ��l1��-7S�Z��@�I�Gs��l�� ��ZwS�S5-Y���i�߭�:2�_�b�01�W��[�e��h�up��P$gTN�|p���]V�֭�9��8#�M�n�V~���%�u�����]���\�ſ��S�sn��5Z^ɺ���e~N�)�n˧�]�ޱx���*��9�_o3hnF���ѿnf�R5%�ٱ��L�H�Q��Z�i�-�tA�gl��zj3r��me�=�Z�9�Ϙ���e��-�{���8|'6��b��y~1G�D��>��\�Ѩ�����{��o
���n�b��'���p�n`�HodO�t�Y��#n���Vkvrl~� y�Ĉ�}w@��ss��,b�8�{K�
�;�|Ym+�xJrM�㠼�bj�;(g)l��O�v�\%8�h�T�6�|h��4B��,�u33`	FL��6/i0��2�T�����pn�2C������ǋ�Hu�������&Y@Ȝ�}�Y8O��t���UaS��O���K����),�k�ky~�i0[#71��n ��]Np�D&c搿^��vS`��S>�Z�Q��ŁfI�8Cm\]��` g��8v#'�ݜ�nθ��ƪ�K���-Ԥ��T&�nÀI�+R��#�Hf���h�qj\z8��ԭ��M���n�Nε_w3��1��r��ೃ�QiX|`�Jh2����F�W�9� Ñ������:�����ͯI^#���.��`�fHVRoh�^��t���>���D�M��u��Ͳ���"2j�F�g݁����,����b�6�T���!�������ļl�'�Mes�����Aĩ�Z�:1��I��`h�L+Q��x,�	���u��Կ�N?1��U���tg�����@M�n&b]6�ʀ!s���I�sC��yn7�xE���� T�~y�$�a�0!0c�
_+3pVc���Mr�%4��=1�2@�������Q6�����nh�e��I�^��|ʁY���F���cf�/�j6��pRBE�/�NL8��0�M\�)<�����g���	���Ԋ�_Ժ(�2�&������p��3k%g�o����Y�C@*z�����*/LKv���Iԩ����2S�ʽi��}"���e[x�,e3d�d��̺\󭖀�|^�f!Z�`'��}[U6[,���41a�Ss!��j��G�#�fX@٬�F�ĸ��Y��U7ӬZ6���M�Гur�<�v�`FM�j�͌p���r�����_j�]wPS�`�Kҷ�Y�5_���Y�Z���͊�Y.)�'��w[�����:���It�Nr3����l��Y!������j+��Ę9폮ZgF�:�y��(F�E�l��jv�
|���`���Q5�S���vҲE�fi.����Lx��>��*���5}�6��q}WNu�J���J&�^k��K��@Ee���O�p��$��cA"�.dn��"�s�y�۔d�Z8C녍L֦�01�~i��*&r]N��r.�"]�hB�.V51�;{�}1�21��jd���}]Մ�nн��|�G�˄>��9��1S��6�fa4��s�����Z���ɥ&g]����2��*�{���WءD���Hu3ۛ3Z%}�Rw�<\�-Z6�T�}A������,pp�x��ӿ�f�D��#�)��v�����&Y@^�.`C�d������$G�B�fqo�JdV�35�J�ʮ35�-6�����>l%��G��*d��H݊���ד�@b�.����&[!g�E9(ȩ@1�,��u�$���̬�J���V�����Wg9,��Iٻ�e�f%�:#3.��W1�&���#B̻�56b*.V�v���f���n}ըY�e���O���U3m��%�_������m���M�¢;�'�t8^����
�p6�,͘9�-��]�����bC&b�R���r�k���_٥�f!��.n�e��ݱ�O����C���(b��{����u�c�۸��q����S�|l��6C�D�{�Z�v�?M��C�Yg1�.�^���j����T������8�T���B(�i&��#�x8�7h���ܽ�Fͺ���֛sh\fdR*G�[zWc	�ܶ�3F����,��M�[���ǋ91Fo@��[sV4�v6�Z>��'%����Xa�,N׭�i���'f�n)�6��d�Rl�As�f�16���0Zų@΅���}���B.�J�?4��:���ZUm=6<��	K��?��@�&��heh�g�bK�N���,�*�Y0jN0�TZw`$����rn��㢟��2�Q)J�
}��"�LZ6g�쯃1`P�ln�.������!���u�xb��e@`s6��)������ј).c˝
S�
���6�Rr�$}�R����h1��f�^�n-����8>���f䘉1��]^��L1:�.���<�l�4G��|v3p���#&��C����Q��J�́9�ވFL�����ϋ6�bc\?�.�j.pNȃ��!�0X��%�;t��X�`�z,��6aJ~4]�7�LM}\�u:����.p��&���lf�1�"n�Đb3K}����Z�Y�aK2qt�,��,fw�e�.����-٫��9`��V��3�M��"N�@mJ*H�<a��2���?�u�Yr�b�dS�Σ��+s�Y6f�k+�t���E|>6���p�`K�$l�R��Š��`���$E^�Ѽ�.s4hB����!�Ͱ��d6`���YX�ȩ �
��p�$��f�Y��u4U�s�J��aVL�N�2[�d�\���{� o⟘�"�����M�6qF��ޝ꾛�e��7,&�y��Jv8�뚞r{p���ևɅk��h&:��0|}b���~a���� <MW�F�9��6j*�� 9r�,ۃ�cw��]����ҁ��|������YW7�Rw�_���I�~-%7�4����j�Ā��rN��"�u�s��ܘ�{���J�uw�����eN@��wr-f1��[!n���+&<�����I1h*C#�e����Yn�UMxү�z.��?��WyX=/R\F+;�ٜ�G�3IaėmO��se��c��?��\3`Z%1��*\�e�׺܎c[���i���_�M��{ݑw�l�Z`�D�K�<��AsB����r6�n���:Ժ��9df�2�&Q��]���3T�:5Ǯ7�w�O�]�S}�d��w������$�;�G�G�,U�e��O�}k�=���zshYA�Cl7%[.�ժ��?SI�ـ��².�t�D�`��5��	��nh}����u�?4f����n~��ؠYk����~��c�����|�^�7��M�D����F�MT������Uc��m}0y��6�x3��{��f"֥�sB�Ϻ�A��l�Q�l��Z��f�+��qۤ��l��F�3s���u��5Kd4}�
6�q1�E��j�O�S~��9�K�Ǹ6f6U@T'D��%�_�0�r������K�p5���nk7��jcd����@���l�6�i���&���7	��l|�EV)T�v��ጄ�:5l�e	���"ef�'���`үVE��"����:"���][4rЬ9�z�	��ew\�YhF6I�E�+�NLX�����[
f��$�+�oa/�Ώ(~��+�|9x����n�ф���=��T0"ug5��}0I��\�˞�U�h����%|�Z8l�k� ���_�g2n��`�$���[^�㴂����y4멦Uec&L���/7K��ӪX'f��_rĄ�n�l27{Kn��E����5����+ɘ	�:2�1�Z���&\uh��·�h三1^Κ�Q�7�r�n9-���b0huh��4pN�իԏP��~S�>�����gĩp`\�U��q1�Q�f��L���C�)�fy���!x|]t٣ ,̐e�LB������ g��v0bܐzoM�52wa�K��@M���M/�j�s��.����ĺ:	�6u�o�J��8�_�f��$��z��u9�Zl���^�l�lQ�I"��a��od��X������s�
N����������\^�d�܋SN��'ȲZH6M�[��hଣ�����-g�ע��!s�<��%�H`X�`�91E��W� /a0I2���킺�/̮C�^'������p�j7'�pXJ"�� �֒?�X��xU��a��0%_K�+�]u��MY�+`����[�'�FV��V�>��7��(J�+���UVs�nG�{��,ՠY
I��,-4G��u0�3u��̸YX�X�1j�����}��!�.��6p��sƄ'���U�H似���%}�h�$�	L�G1����91�Twh����4�����j)/>1f�n7S������}w�Bs��S�_�S�0����\8�t�A�t#�кު��U��Φ��,���Y�C�2�I���r�0
�݈��9ƀ��Z6� 9��j/��qA%�����G:1h����"Pہ�
�/O�dQ�}����s�m���AS�.��݊��^1S�:L5#��#e��v�Y�Ckj��0�Y�C6յ������36Yw�F�[妒���sƪ$5��9B���Y���㰜K�&�nY.�uT��M��BdcF�0�LR�UYV�m�����x���K��}=x������}%�&j]��]K���/N5aJ��3��l|e�BO�E&I�E G�j,hp�d�^䥿��O
i�߸"��M�����p&w2=6f�O�����}Y�d�Tv�����]fI8�Rw�_rX8ZbԊRw�����8�$2��-�EFN�&�Q#LЬ��/�6����)� z?��6I�lΪ[�I�f�m`��?ǭ�m.��?�����l*�O9Tr�ȉ�������jVC�暯�741�ʹ�ظs æ�&町y%I�9Tj䬊����c`y�9��$��j뵩;�L��n�+�DҲ�]���P���D������7�~j�)�f̨���l@La���pȐA�T/R�6�_f���(ur��-��\M2����3�A7rں�Ͳ&3�b���Z�ᳪB�z��B fa��1�=��������C�F���0&���*j̐)`qT���m�L���e�@K�R��x`{r5`�$Y��o�n��S�ج�C,�75k��7l�21�_6�����������[�5~1ۡ�X� ���QsW�)�rR-Z3��Zg�·hx�7����T@�ug���l",�-+5��]�I� 9Sr/����Ǟ���������-�M�as<��A�ɲ(���X����O�}41���d�\3�D�֡9MȌ�q�h��g��V+q�yq����Pc���&��uO�J�x��ĥ�`���p�����s�W�5�ʲ_�T6�t��`55�+����+/5b����)�.���8��s�M���i��qcFN����"Pہ�
�/O�dA�f����3���o��6���f*W���L	~�O��4��˹��N4dZ�.���F�j�j��n��>;��S��7�.�/��p�.)1h�a�ss�΁�N{�Wfa��FhR�^w�69@���D���-��ZW7aJ��X]��őP�6�fX�I0p�ɯ�6+��+�-��������Ne0`̬�i��%jݓˑs_W�L2�0hȘy56��r�4 ��9f�c��n��P��ɽ�w�Zy1����O�uP�&����(C�h�;9n�mI�xk*fݶ_a-;��h��2;�$����̒[^dڲ��(ss����]��=�ؤ�G�s��J�[9ۧ������E/���U]Vb�kC�g�����Wᒻ9�m�M��l�\�3TMM�.e�A`���30L�e���������ԇ?51ub��f܈)V�Yj���N�Wa!��˳���x�7>�gߦ�����b�fS'�2�%5`Sw���+d]W�r��`i�d"6T��"��s���~s���z��
��_�sn�_D21B�4�Q	�p+Z]N�f���:���&L��,�����!SݿR�R�vaS�9r�<�
:�'��Tg�P��<'矛SyW���Zfv�+�&ƺ��w�1k�&d�S'Fh���l
�Ѡ9&VyM�)F53�t<�AS�x�e�D��N���9G�8��|�lκ���ŰzU��(�}����Ĺ_��F�!j"��e��e��$�s��x@7�zf�,0p�
�V��b����B,簸�fV��6���O��Qcf[2W�FD��.����,�#�.`N�͛.�9 F��!�MwE���� T�~y�$����fu���虍�`��ڴ���96d7��
1S�bsb�WQ�1s����Y�$��c l��i���nW3�@S�f�L�h]W��%�f���2���5����u�T�qn�܆u��)Ćs$\14����ٲz�iy��u�X1��6lbXt��9P�1s� |�\������(u�νY�-�#�-Ƴ�ǘ���w�͠�u�d�p��#Y���|COn0p"�e��{��ld�o�&L�W���ΊU4ݵñ�����.YG�ʢY���}e���r�M�͜�d����W(����h�Ĕ��y3l�T�����`��DW���*5p�պ-h.6ɲG�gw�L��J���1r.�3�d�S�[�r_���,�hU%-�ۨf�h0W]��t�%�|�$]ds�,��|
��m�r�&3I�#ՁY�ۮ����Q��X���P�&]�2��:���)�@nq�����p�Tȑc��_�15��"�DC�L�[�C�:�iU�3ln �f�*/��g����8���?�.; ���� ���1thr��U���u�8!�(A� ��I5'H`��9��23�sc�Ԧ��fc+L���Y̒6S��dC��QXq�^�fq�!������, K�M�;Fn����if(��h�������#g��I���yL]<4rjb9Y�f��$�"��P1b�T6n�n�Hmf�ĒvsM�Ĥ^>KA͉qu��X��b����z!�����BMX��R��l�Uj�ȁ�T��d`��v��x���trj�K���z���T�����CFN��Q��z5�]���I�� �6���BՑ�֏v�$ӣYx�1��5b*��|�ؚoN2���-�۷�ٸ	y�h�ﺁ��j�j�kv���$_Ճզ��i�e����M'	��~�E���"��N��u;cT[Ю�s5�t�q�W�P�&Y��z'⡤�N�uz�����a�R�9P��u��F*�M�N�Rv30}�D,Kq�=<���lԀY��s�tق2�Yo1ߒe�g=�䬐������*E)�����rV���Q��l����:I�%��C�XM%ͅ$fr��&7��-�����>\��[�kq^ȉQ+B����\�W'�<�7a�j�)Tn#_�5�ˁ�
`���d&j]&Ѻ�۬�����%�������Dk&�N��¥��!5��L̓�������Ksɫ��M"3���Z̢:c�����T0�P���l�T�ٱ�&<�#q�=��>�,?��m�>;���u�fA�Hn�� (��b��k� ��X~7z���:6HG?5������F-b]��`.,2��2aJ�f�h6��KN��sO�d�Vg�������sP]���E���z��I������a�6n�T���fV�`x��c�1�Ɩ��u	�oz٩93��	O�H�#3 �T�l~��u�8!�(A� ��I֦� �.+��-�l�K&��g�.��V�п�Q�L�}ͬ�&��AS!K�-]�b��Ͳ1��́��v����uU�,e9jܠ	S��y�=�#&	�h��N5j6f����sQ�ᇍ�$�n�k�5-���&w�Bb�dt÷&s$�ٖIw��1�z������b���f��=֗�J,�
�+@��]�d�Q81ew�|]��M���lv�hԄ��huQiFM2r�����Y�ۨ�]�����G���kg�2h#ㆍ�P��'s��1#')�8��Yp�ܑ�T���d�=�+�f]�P�ޢ�I��������Z�f+4�2��I��v�as.�����Ψ+}�o<�n���'B4b"�e�<�dῡd|g�;�oh�k3灘0Չ9�V8�$	�Q�����P&ƿ�_��0[U��3'c�+��-es����T�Ѳ�Ӡ��~�ܾ��Mĺ�S���l6��
N�ӣY�͕�sd��H<��13��$-F9���csH���ZJ��͙��[&�r�������D�`�AɺG@���r��۲1�鷏a�Q�Fr��rn����� N�Ll������&?�g����0}uݸ�v�Z��Bz2$-[@��	x{Ԩ�X����YJ�po�L�ү��3�܋�>���F��8���V�9���6�&���-�#ƍ5nਉ����k�fu[����5h���
��$�>�R�:֖�u_PЄ)=�#�T=����׍ͭD��\��=<�%�~'k�;L<�����k���]�'4�j<�{� ,��&�~��l�np�p2�=���Ҋ8!�(A� ��I3w�0\�8����j�@��6݁��9Ю�
:؛�����M{K5h��7��\���Հs�"ud�Qy���I�İy��6ؐDF�i�f�J6	�Ġ�04g|q��zM�`�p��_�._��D�����rY���N�҃9y��e\a��z�:�VCL�E�s[nĺ�1���o�� æ$_̬�Ҙ�d��^ͽ==�/<n�Y�r��D�*���7��ɜfԄ)�9�r�!0�n^�9#�0աY��1r����/B�y�K�*�x�:67���M�>3!RG油�r�;a�[��/���M����$1�D��Lx�J�I���fۛlf����L�G��dz7�>WLNQ+�,��b8���dQ��r�±rn-�,,2��8�+Lu'4nN1d��k��h\/2f���(u��ͦ��`�� J�23ǫ8�]��vD 9���?���h��IZ��Z2n��U�u[�++'G5������z�:Eڲ;ߞw��)&<{;7/���Ð���Yw����Es���Ӎ�0Ց90�q�)4b����.:��l�*�yW8��"Pہ�
�/O�d1s+� �e�Ac������*k^��/����o��f-'�.��z�h��!#�];������������s��Y/7[�Hݦ��y�Rs��u��|������La
G/[7kz�T��n�o��u��$����B�f��C����l�����7�FLx��ܭ�4�J��i�YbĴei����o�r;��^�`�z]��)�/�f�s�1i�]$�lﭙ�"L��0s�/�08{Z5j�#9�I.�9��YV������7�&Lu�I�f��1	���EE�X�,^�r��LX�*Zݕ��%8�Ф��n�lN:6qB�f���n�28g�kVZ��d��<�q��:5S��Q����L�^n�:9ǒ3�R������7�N�һ��pC
�.42�p�291�E�;���@&ƿuх&G�`r)\6a�{��e�f�,�qHQ��s2��۴�$H�Y������9��J%�Z�E��.,+��Z��`��r�Q�L�<���U�YX�g�b~��b	�VA��e���IL�ң���������7��C�1a�3ܸA����/B]�-gI~�{r��)E���� T�~y�$k]/E`�,0h���Sc�6�����ZQ6r6��+@��3M�b}�iَ��|1��MµMm|M�8M�0խ����]AӢ`f�ߔ��r��[(��:�1&�Vo��6�؄ɿ�/�͊��SA���M4p�L�D�ͮ�R9Tmo&<|[�b��݆3�����Y�F����ԩq�L7�Z9hĄ'�K6�� �Q&������"�jbB�j��[��Α�ۡ���oN���KQ��یf��s�oz��	��Q���Y<r�^Bɺ��as;ܸ�oif%�2�����p��=+�n��9����4l����7c�7g����l�r��e�&Yw��p�OH4M3d����,�CU�71'�Q��5u��|G��
#S���c���WLT>F�����aY�	#�TEg��A#��>Ԇ	�Q�3�B^jf��Kᄇ���*�#�M&<�\C6dV��Þ�aad���\��-���D&<�\J�g3�C&<\�Ճsn���A�q+�E�g��F���⥸	7�0��uA��͡�3�Rws�^��9<uॿ�K��%��th.\2������7s
�F�n�n����rv����@3IBD1~e6�t�L�d�
R�lrn����³�zk��Ӻ�+�cf%͐�m}���$q%�A�.����H��T���re�E��廸O���50�!�к�a��f���o{^N�a���,���^G¥^4������|'�6�f��Ik���Q�AC̢ObYmr��zqS�܀���f1&���5�c#�`X�l^��s�M��ԙy���k��/J�3p���8c����kYU[9�4�4ɺElf2�Y�ՈX��[%7`��Ó\��'g�(��ġz�YJ�+�̍����j��|�ܓ�Q��q��{H��d��p���4j�.o�0����68" 1I��I��Ϝ.Ssbl�FͰ-��`)�Ȉi���]�����9��"?6ѪR�C��4aH{8��*jG爛*��s�3soФn�s�-�;"��հ���d&?bݣo�bln��v�:2[o�
�'�/���l�U�23�`��Ǡk8�.Fΰ�B�G�1���k6k�fu��N�n��6�z1�:���rfl �s����M��3���_����D:j���6�xU�_�:E���� T�~y�$�z�S`�w�u��D.h۠�MK��V�1c���7S�߮�*�AS����Y��)���_�]6��P���B+�������v٠9����#3N�Q�wI�W^̅~�un�Zbj����L��'��c��˴�WzYb�V̐z5����e��@0Kf,+�GO?5�2j̸��[�cia;/R�E�[x�,�'�Q��v���s]6u֞P���|���f*�����c��.�76j�:�Yޭ����-@G�Fbdw���M%y|Yʩ�s�V�j���4h�k�`�2���M>��g�*@����²�&�ש�^W�H����u|ޫ�T�=��Ǧ�eSe^a��o�d����V����K}|�����<ݐY�jե<�ϔ�;i��g3}k��w���.��$��sv�,.a4p"�e��i7vM�ҳa��`�n̸��?��;����D�sޛ1��I�M���zb���	8jb�۔�C3l������5k('�Dr�0�s���e)���Bj��9P�'�@$�e�Lݜ�Ro������/����=�Zg�ޭ��;�$�/��Æ�`K��j���^��h��$ӣ�sڝ�+g���������8!�(A� ��I�)�0'�ko��G_�˹6��x��L_�ֲ�>p�9T�ըi-ljӇ��&���od���7"u+\��]�{��s�fY,{�.;��e��&!��Akp8 S�,/������6����}]�D�˾-���'1aJ��\��x����ﰸ�bĈI�hՎ.2"���	��j6��.�󌌚�"9Wr=�e1Ư����^��W����M�9?İ�j]�́t�fV\8aJ���	��{�V�9x�Y�rܬs�"�-T'��MlvCI�"�-�-��J�j�$�V���F�q�x؄H]C�%�ً+Lu�pxc#47���?�28g�k�?	�j����lQ�6����#N�ܜWV�ʓ�X������8�I��K����r�d���w+h���Q�N(8h"6bАI��.��ؠY�cu�p�T��@ݶn���M��@�RfN���b �ꝟn<1�Cn�ŵYpb�R#F��_��H���Y9�|�ZSN�Sta�Y�+�f!\�����K�,�M�����p�¹���ɀdf�,K���FL��Ȁ9�ݠA�f)���.:�ݬ/��*SN)��v�����&Y@F�}��֙�´vd��i9kȦ6XVs���c�uf&�.ǰ��]�Ր��4���q1)��}����sU�����~5���l �c����]&h�n�Ú���Rʲ�nioh�?��u�f=�t������[3���,[ϕ��'��W�N�b�V�d�XW�_6n���8d���##GMq��w��fR���`|_�26U=8G�x
���6����p�	����fIk�%ҟ���q�fm�L��`6����ԁ�M�������V��qQ���HĚ9'�e�]��F���8nF�D�J$G����uk����[�E���?8/.1Ux����;���S��;�Ĝ5�Jl|���1Կ���L��L��sZ��ͯ��d�%����Y��Ux7�>�Ñ�L�j�ys���d���#�0�&����M��ދX�	~�Ǯw�	S��y׏05øj�18�y�dz6�ځ�|���9.0n���Q���J�9�Є)�;( �ܞ$��\-1,6#�hk��k�&)��lĘ�X��~A����O��t��p.U���=.�g,�+��v�����&Y@���>�����k9r��aS���
Cf���n� 1S�$fI�qsU���*�5�f٭����Q�V��=3���$�Yp�eu�,5ၤScVc)�yWX@�~�ٿE7�I�`��O���LF.8��-Ԙ	O�V�!2t6l�$�7J��s��&�[�{�����4�T'� ��N��p^�����r�ݧ%�f�O���rk���D�+�ofcj����m~�/;8r3'Oŭ�۱y6�.�DY/�r�`,n�t%��и�5�@�uh>p���(u`�%���6N&��c��9��Y�0��.��µ�b�	�fx}}�	���7�Y�KM�M� ��tS-C���o��Ib&��(ur<nֆ��IZ��.��-�BcgMVQ��8��ܞ~A��G��Ư�1����#�Lx�G�7��ـ9T�:E����'L��TM~����rE�9�ڴ���Y��ê�Y-7dR2����mV���?�Z�n�����T4\��=_��^�p"֑)u�g.��FS��8�I"�u��%�Zj̸�p���=<�ͰI���m1��y|�A��ek��8&sHOԽ���æ֙9 -7��p��C����<b^����R�Æ`�L��Y���Sa�u1n�11ug+6��]6�{��e���S���B^.h
���l�����'���F6��S�̭\TI×ڍ�5`��&�	N�|[��$�b9��[�����M�X�E�;��d�/;1b�'�SS�7�^pl�bb�~ƑYPʍ�Zw��9D�Y��$�C�f�l�q�ɠ�ꝏ��X�d��^�5��*��e�[��z��34I���j��e��4��y��zm7�۹rb��p�TR��K{{��un�i�����������r��O����r_�fj�sdu��q�PM���xz�D��B�PAha绘�� T�~y�$���!�|gsK���2`S�V��vL/Y1���h��cs ?��QC� ���z���6�F�u������N'D��2��-����O�J40�~���6rРI����:-lf�L�$�7��'�i"u���|Q�F����Mp#�G�59�m��B.&��gf0�nj֥��+d;3f�$Ql����Ő�~r"����ʽ���	K�%x1/�!M��C������YL�����_X���{�,v1b�4��P��n����i�d�PG��̨Q3` '	@K���K��H�TXޖ�B��Ր��͙�fџ�k��Ѵ`��y�s�ƨGf#k��լws�3��[�s3)��x�=��7b]&�E [�Ef&<���Y�@��n�T�d9���m�s��%�F�hV���Kͅ��ŰI��`����Ӥz�:�YٛfFL�_�,Vqy�Y8j��Ku�n`��u+��$P3�!Sӯ�*,�<9�j-��E��������h���ą�(8�#Ve������!w݄'�}A�,��Xm�v��"4�9I�TwJo��F#I��ԭ�)}&_��4i�5�����
+/F�fo�vq�us�6�d����u��峐�y02f��	Sz1K��s��T�Ϗ{H=����W~e�1�Z�It#&��(u���^�xzk�"N�@mJ*H�<a���+� ��Ks�b4dθ��W�e,��ǧ�%b�so����T����9��I�-J���/��\Ұ��
�,g�,�@�.r�A�^GV8@�ub��Y@5d�iI�����hb*�6��p�}4[$@&Z�
^y1dJ5lذ���/J�%8���!3|M�_�h���c���J�ՓƛYo6��f��x8�_�ۭ3�8�F��QOLĺ���/�����}8ҟsKQ�58��!S�_�5l���dY�/9�k�vj�R��ꭜ����M��&6���;~nG��й��hF��R���f�RZ���-l�+�dФu���9=Ȁ)���^��~v�O�0�'���l�~/˪��AЩ�Z�:1jV�$Af�I��N΀���XK�?p�������U^ō��3j�_�uX)7dĨ�X���l��md),O2�H�c��Z�W�M1\'D��%�_�0�g���#�z���8����Ԧ��-_v�����c���f�޲�7ef��Z���u1s�2���h��J���P���o���.�D]�b�Ą�̊�Y�Ȉ��Sx�{���Ѕ��	���$����Z�_f܄��pQ�87��M�@5\���Q�6k�Tܤ�G����V̡g��D�z����:p��n�K}��ʁ�M�:1�nݖ������5���\�����|���a�Lȱ��gCƌ��4b�T���A��M�I��n�jVi�u[	7I����bn�ԭǖ�b\�?Y�Tϸ����;�� �o+'���|M��Y7]w�S�`�N�o�>�^�OU˖�f��!���u1��>`w�iy��9)��o��F��0V�-t�_���3�$ӯ�z�ҹ�Lu}��̧�}1��U7�R5A����m�^&���;��\��Q�j��u�[��I��,ī��VdWLx�e��Һ��$�^�� ���\�u@S]_��C���	������f�,-9�Y4j��Z���F����f跹�p�d�3-��anu�V\8��D��.=�-��1�.���Y��VJ��(�UKLʖ�*�`z1�9#����*�	W�a��X�����u�ू�B�(�G�;�9�az_�,���6�n�cA#�!��9���ɯ��-�5\91r��0�R���}{3�9F�Hu���附�΢�� S�ތ���S2��55�{������He�8!�(A� ��I���0'� .����t�k��
�B%��*�Y)2@���+zv�������%�0�$1�%4\����A������J�ѹ�l�E�/Z]�Ԅ�awmC�i�� V��قfq/Υ��ed��j�g�5Sq��bN88�a���l}�����\	�q_W��L��uK���`s4���b4nn��#�m�Fͺ-��Mxү׭�i�.�~y��5l���7]���\%3`�)������B��� ���sHY�+H�2s�b�ud3/]8b�D�+�2�e$1����-9ر���s��-�s0<u�E��w���E�C���j�ιsy�X��:�:2��*�a3TN�?��Zf�TփY&'�:]���h�,Z9�a�d�����{y���l�,�wx�#�|�꼖L�3w�]
d�T%��>5�02I�F(;���_�m�*�?Q�Z�v�Prc��7#'�ȳvS�j6o'����Cf��7O�Q��D�u`��W��Ҍ#��s�/y���d6rя�
yѓ�Y�U?m7��j����s�'^s3�oA<�>U��Z`B{fЄ��y�14hbX�n1�.�{*&������[n6�`.��v��j��n6���j����jC��Z��e����-�L���܌v����2Y���>�ɥ?'��M�����.��QXR�9D�fd
�漢�C�����и���Ɂ����������Q�pp;7�`�9z*���Vl��!�Y9fb�;^�#�_�Ds��l�� _��Gᛛ���bN������"�Sȼ��9�7i��VŖ�9���l4��5]�C8j�\W���5��X�z�ZI9F�.��e��9b܄'����j���� ����+gL�yl��Tg�͐�̡�MN7��5^R۴�l��-�lI&�.�k�"h��D�K�t�+�H`�)}��8"�5ؚM��"N�@mJ*H�<a��2�.+�`lZ23p�,$˩6�Y��t��Yn����"]Fp�vM��Ȩ9�-�k�&	pQ�%9jVd.!7I�ϣ�X>�af9�	�:7�6�*8n�u���m�`
Ŭ�����\����́kd;)W�S��$�����>T�����2b��I������nbXu$�����{�z�d���Aӡq)��"�N�&`�,`�2;S�u�������������a�.�v'Wh��4�7j%7���QS�������P�M��~k}'o$���jV���I2u�~�lFN
��	��Aҹ�h�R%F�!��E���L��ۭfMʏI��V���M%�/Tl6�f�˛ż�k�$���MC!9+w���& ~�Y*l��5��겱jN�uy$8��������:/����Zǣ�Hq�N�#�a3�Sc&�_��es,�9շ���q�60lĠa�e�rX)3h�q�oY��^y9hz����,7)_��dVy!uc�$�/K9u"/�mw�	O�U=�ΰEA�L�̜Sf�7ɺ5����Z����������B�N�1��D��a��{0W7������d��⟜ebf���1$Z5n���_��z�9^b�VͺbV�&_�5����c,;��fnV��&��%�F���9NX���d�V��G��gs���h�\($��b*���Y![/��P9B�△��9԰I�Q�:3�^�9j���6�f/�#9�ަ������<�T�x�NQ�R�Y��Y�Z��$�i��V	Kf�������6jЬ��vֺ��Q��a%�Z�Bg�Y�����/V1A6w�&�~�Y���Z7�����1T�qBj;P�PA��	�, ��0\����j{eѠ�Mwdcd��U���r4S/���{5�.'����ZF�7	����G:@!R�+g0�`u1u`��bΪ�R���`8��`�&QźhuQ��r-�M��Z܇Ik3+��ܨq��jw(���kaZ ݰI�4�qub�RFͦn1�u&���H���.:���f~��|[a�s�`�Y���}J�Y5pVN�4�PvQ�,m9g9`����YhW�n�k���Z.r��`�Y"��\j��ZVOv`�_��$�n�U��EW�.���,�nF��$���g�К�#���Z�0�-\�q�f�쑓�-J]tF.���F�'4��Ĩ1��%�&Lehn�"<�帉�w����^�"fMݶky�_M��{}r�����R��Y��,Ր��&L��,�3D��9��[*���b�V2a���r�dVj�1�����#?�Pm�LB�
}��q4©�#��� �t��ashg�L��6(g1��:-����zN3��*I���!l!#Cf���u���F�l218�f�����j��p��`�4�H���c	�9yݸ�XW���Y~�nhԄ)����W��dS�_�� ����Y���o��ʪ[s�N��I��ln��RS���z���0C&�~�߇�tQ���e���,0Ir���+F��K�u��Ƞ9��ȉ��������~]�}sl��r$��98�]91�$�&b]J�3lY��k�&<�KG�%s`������� �8ɲ�lYh�3U���F�@���UQ���9tG��M���w~�7�&�73�s�1����}3��wݴ�Z\����e~��!!X�b*t�!�i�F��v�����^P����P;
X�y��^s6d��E�͠Y
�/6C����= ������n�r%nz�un.�����ʿ��,�5��M��zʇ޾�5P�.G�G"1hΊ��&ZY
8�
�:�RZ̑b�XAsR�G̦�Āɝ]�wn�@Ժ����YP��`e�ܴ�w�r�DWI'D��%�_�0���}�Y�V�����D�۠�M��n��/����G�e���p.0f��7��l�I��8^�͙Z�]y7�xT�̦b��u]�'�r��p��X��Ϻ�Q���YNnj�y^�k�&�����pn�Nr�\W��9hVz�b�n,Y�nN��ۚ��m��O\z6�R�#����'�[N]�Ȁ9�ԄR^g� pK�����?|.�%�fI�)�1sR.���{���ི[�!S�csz/F7j�B[�h�ذY���4fV�w�K���e� .�Զn2�� ����);ـ�f�.�N���ݗ\٣)�V�:5[����K�;u��y�����[#0I�����1���*]t �k�>j�$�z�¥���&\u�z%��]}:�W�
��j�.��15�U�ܜ�8��9��H�����/�5��74I���9��OPU:]���8��P���'��gס1��w��^2�8l��[7jJٝ3��c�fo���e9�I�Vb��D�� �~j�r�>��ҥ}F�!CM�Vĺŵ�ml��DL
���Y&�26`�^M2�i�n�gUH��K=qB�21���s�����^�ߵ�@R-8�t�/1�u8b8��Ϻ,u7#ة3s�[��-
21�ZA�֊yd�T�X86+�����ׇ����Zwf���K[N:"��74n@���`� ���\�[G� a+61�9�����e	Ҙ�s..���0%?������Ժ���l�*9b��O�5#��.7�26����3�E�eu�?؅�-4��-w3l�T������j�H��2�����]���Y�N81��ȍ��c�j؈��^�e�F���M	��ݟC�-4f�ct��g�r[��eS��Y�+T7/��[��cs���q?J��R�����Q���#f��15�����Ș!�,���l�������Is݈
�K@�4kx悉��g�Zo΂.�v��tZ�1sJlW\W�	��@	B�'L���� s�����9E�۠�Ml�V3��u1S����9�Uh�k߯�r@SA�hg�v���<w��ʪq��.�I�H̢13Z�)�_��t��A�0��>`��QS�^��Y�p6�&)ۡ~�����"ZY�mI.��P�؄'�1i�,��),��ú���L���r�M����6��$�#��yd0fV�$�����ȹ��7���{>�qN!���ΘQ�:f�d�򮃹p��Ⱦ,��j�A7����'��ԨIr�̵:���0j*���eqk�?�~�Z���f���M׉As b�.2S��ͪ����f���y�/�uj�< �e�@I�#չ9D,%5�I�7�$7xMհAS�_�eu\�!�&Ʋ��b��Uh��WaY�hG371����t�\�u)˗�a��^��I��f����fV ����p�VS��ǂt�W��s���3(�j6r̮Ժ��cCf����A�3ߦV3Eh+��N�e&k'�I�:5�.�ɲ���&kp��17��>¹�l�$��cf�.�c���23ùe��6��c�xٚ���u9���%��P2aJ������Yi9����8/la�[ �ȹ2��О�/R����J�!럘��/e2pj�3힨ac�*���q0U�#h�f���S'����W8Ex+ ��,��F��Y0`&PS��a�_	'i���]�w;2��ͬ�FO����ʹEK���ٕR3L �~����+����M����`dݏ���k(g`�͘�n��9W��?Ӓup�΅���W��wlޯ@:�����r"�e~/�����pC&L����ת�u�1sPZ�#��)��v�����&Y@̼�0\Ε�=���t^�۠�M7~cdجȪ�y̵������\	9��m�.- '��'ɻ�p�8g�8�c�L�`�LC�6�����K2v�Va\�u[i3�X1���Ez^&�^o;����Zv�W��J$|;I��j�
"k$�� $Y4`�����\�_�Nbb #Bْ��ٲuc&��m�l>E>Ƥ>��,���U���3�>:̘I2r�O�۵��uĺ��z-��	�7h~٭��0S�9�l�W'Y'�[�E~�;��?�5���8�n��XzM�Ժ�fe-��O�-��8;ᬭ����|Y��p����Xǫs�t��,���.�lb���j�ۡil��]�fuŘI�{����%�<�D��r�-�jS����Es�N���ʷB6������I��Vv�>�=3�+h��S6�H��nE�l�bo�'�v�:2�0�,35nbЄ��ߎ#�ME�&��:��d�=;$��(n*��1s���SpE��8�n	�����>Kl�䜊���Y��wc+f�M(�5fs<o`�j�t��lnG�у�����E�&z�"N�@mJ*H�<a�d-ש0\���_�b��v�k�RG�12wrl�D���h��g.6`��wn��r$���-�u}1Ud6��&���I :��9��Y˦ʴ՚-�NM(_�bаi���0D��7=��p9B���7�����	Oz3h.�ps��$ӣ�����]w�����M�8�f
�� C&p�`F-8hN�p@�ٽ^W��z���s���G85�jS/s��[�DZ�:1[��!#'ɉ(u�`��F�K������s�Z�
�`�ܜGSC&�Ƴ���>7�r6��O��:`.��@d̄��۱�����核��M2����\#4Gg��@p�.��o&I�Hu�k,�sp��,B݁�u���j�@w՞� s++���psulb_���M��j��X��c[6l��(`.B�ؐx�h6�o)�AC�W-��b��D�K���3r�uU���}b/\璜�~AamF̷H\��~}����-�d��+�T+B���e3��ed��x9�E��kfF�M���3�����u�Ӻ�c���jV����к9�+F���#dY�a�2�NR�r^C8p��ݨm�^��֢Y/6��f��.�g��uX;5�+�0�
�Q3��AS�_�k&�3�̌g�=n2�oQ�,�hSp���K��y6n��f��1d�A�_��E�A3,"�e����[��Ey�S�(;k���.��(�r2d�l5H8Uh�
G� �Q3�,����'��,�8���5�3P���l�ĩ�n���{ܺ�X�`��Ĩ��)��N̕��fj�s@��l̶᩻��ʦլxץ��PwH?>��A>��d�G�k��lΌ�U�_���y���m�D�K��Pg�İ	S�(�KΉ�~fj�"N�@mJ*H�<a��i1@��0�M�6b�.2b*[��"mlE�l|ŷY,fj�n���m���q��b��Ͳ1������!R��܈sf�Q�M��;8h�8�~���wm�PTr�Y��ۘ9����d���+�g�.c3�ܙ�Mҷ�?���Jm�^�]9<g����&����G�7&���l؅S�1G���MSa0��C½����0rMB����[�`�����O��Vr�FμՁ*u�d�X9�7).��-K5KP�eS�z��b\�h�TX~Ѻ-��s�u�Y*k7d��Ѭ��������r>0_ЗT��;î��/�ML��m��_�J�u����Q�Fl~����_�l�T�mz���0u��	Sݥ>@��f�NBu��͐Y9pF pb�;���9��	N%Ȳvs���h��[o8#�i��3�l�͚�hb��^�w��X�rn�K���laJX:�؀���n0�3��$P��*�Y��X�
j�\Xnݡ@N�� o��m ���y��������Y�܀���y<0O�}����ͽ=���`�lMV�0(�n���j�T��s�,�7gC1V���Z�e�\�T��u�fݗg�UϿ
r��Z��X���,�f�wA�������W��nI��x_C���G��X�հI�M��e|�Xn�1в <��+)�l�`�4_b����'g�A�.5'���1aJo�f/��!��B��p�Y~`��q��4���_�_�sbE_nb���lܬ,�ӑ��j8��{�>ԹQ�L�f�]�ʊ�`��1��f
*��v�����&Y@̜C}��&`��V��Ksk����)���B��545j)p��ӄX�ꋗ�	�pk���j-���M���r8/CCf (Y���A	L嶜Ӗ�2S�&�e��3_�E�F2�79�{-I`R8x�0�r�@�D�S�F���YNnب	S���-���^��i7p��1bR��2�9��,"8l�a���l�9�T�V~A��_Af�����	���XPĜ�`̐�j]�o	��P��0�D�k27���c7/4�W���Q�:4`N7��I����:zհI�����׭
-�e��~��<Z��)[��'���M�p���#GM��j޹��������sd�qs�v��)�Ħሁ�7nVc���{6�R��	ͦ�,K8d~#�v��+��B��m�91�E�� �\�l�,�1�E��pl4p�23��!P��ݬ#6�M"��mφ�8ph�� ���S`��)rsl
������l�
��hl�l�bƤ�sZ��4����e��F̆�l`}݄�Sh��Y�e'�,�
�Qӿn]��ЅZHe�A�ܤ�DL����94KQN����uG���}��W8��"Pہ�
�/O�dY�u������-�!kuּ6-8�k�l|��f3S�Y�����q��/^̛G��9g�hm��ԑ���-u0�:Yw�؈��L��ڳY7d�2	Gn؜Xp.���7S�;���2���d��{A cf}а�.���{iF�u?�Ó��@�U�5S��΢Z
bĴu�n�sZ,��HN��?�Ԝ��ZT��as�n��}L���Y���2�q��g�8������d�C���0�����;�TH[>7o�,D�&Lu��p#f�#GLҿuQ�>��6~Ƹ�c&D�>oy	�34)�E�[��7���M����QF�{��M�L�J����]�Լ��
�j��ͣ�'�~�M�y���X�ҋ̦�9�܍��d%�,�����"s��\9rb�:J�	�������.����ӓp��/�0�;Jݲ^�f�l�71�Rv`&#��#31 �f*F�9�p�ͱ�vh�e��g��h���+���d�ey����"+t�.��ղ9�,�E&���,�E��2����p�ȹ�b.<5��f�ܢ%|�|���-���5B���"�E��ن�	xVC&z�"N�@mJ*H�<a������e ��[��j.�AMmZpVw���Km5@����:.76�E�e;�E�&��E����ޅ��U��Y�]�b���Иو�d������xY-�n�vC&Lu�z����h����>L���]*f�ҋ9փ\D.no�u@1&��b����y��NLL�915K|���	Oz5�e�l�\�0��f�==�#��a7�ᑨ$&����t.ԇ4��nԈY:�G���KQ���|�pV�'L"G�##��A|���������Y�+A���\ 	�\]1/�n��&��Ag�O�$kd��mM!�_ץ�O��j,y1l�������3`*��ۮ�pv$�\(؈X9��t�Q�J�̊{�:2á�[56p��/80h�\�/s����(U�ټ���Q�����Q�3h��������0�s�]6��0j�r��р	â�Eg܅��V,�r�	Nx)��f����0��\�U��n�#�1��R����7�R^���&e,.r6�N��j��	����/�ګq�&Lug֡a+8&�����m�s%шi�F�,끮�q�����Y��;�i����m�L�0Q�_�%�fm�N��Ϋ���6�>��M���>�����]��Gfx�Z$�bs�Ȥ����=7<��#�7R]���1tI.��E ��Ŕ�n;7dn����24rl��e]����52���׭�ytլ|s󎮛���i�([6rฑ#g�_h�^���&I�u9#7u�M�@��ܡ4���Ԭ�!m �٧��/]����-黾��4I��ԉYl`V��"&��-��Z�L��h����������Mĺ���<��*9l�*-��L�^u�7����Y1u���b���"�|����Y�E�&��kxPe�fN�Lu#fѨ�)ۄ�ef�,k2����Y������I3 �Rd&������Md��z,�E�~l;�h��1#�b<z��D�J9�d��:�	K�3���R#S�Z<c�_h��ɑ�fɻY�%55��6G����ԁQs��ئ%Iw#��2l���ut��W�9���qT��̔nb��$Ňsv�9��\�r*$�1s������LF�GQ#�˖�!m������ycf�LӉWyY�96Wd#I�<Y�Ρͺֺ�[I7�FL����閆�N'D��%�_�0�2@�.`b�]�bq���ڴԗ��#fl��fj�j�6��W ��7k���-�2%\c���R3��	��[J�͈�o٭���\�c�zǑ��S���u[5G?�dݚ-r8�r(�֭�f���!���2�Sg6�i}�\�	�&�n��7s$����e�H9de�6Q�Jr6�C�9�G뵎bV����Q��(g�����E�[6d�E�=�N�n�I3r�L�4�,�k"��ꢉ�o�/�M-5�q�O��	���ڠ��}�+�&���K9�J�s]՜Dd��)�݌��n0sqr2f�@����q�6����ͅ���l����`�2p�t6�u�.5[�rbX�lWI�t����ʧ�>�Tj�l`�V뵭 ,��g�7[w���B�fUj��\a'*���c�]=��"0Un6� ��|���j��9�����.��
O)͑GL�҃9��,�ki�LuΒ\�6���"�-�r6u]/ 61`�Ό�#č5�Ij�!����QL����g�͗�7�T6�&b]
Hǖ�#�0c&L�ј9Hop�nL���ޢߨ0`b8��dƎ�!S�j5�$�8�Qo9��*m�本ƣ�@��P��dz9Kr�V�����&+��v�����&Y@�:���3��5��4Ѡ�M�¶��Ld8۬35��]0��i8E�e���כLR�� ���dĄF��Ϋ��{�,�?p&�ҐAF�i�T�L%��<hV�P��ǨܽJ�i`�prN�޹	g����f����j܄)���:���3��~:/��M��$K�}A�{e���M�1�`J6(�Resp̜n�8�/��O̲�#&L�9ۗ�}_g8�1~Yb�)��&<�7u*�뉷�*A��
\�rܬsN"���uؘ9r�I��N��^��=��z��:�`Ԑ	�:2���%8�W���3oY	61B�8r6v�S����Yi5I�<�28#��Tt��6�G���94-K9f.�u9�*'�v�&L�ѸslRL�؅v�!�JN�uQ�n=��,�b�l��� 49k.fy��'\|�P�����{t��(e�o-�f���@�fǢ��V��1!g�T1�mj�^2��\���u���䬖�D�a�*����B��B[�M=������pJ����٘�An�Z��rg����o��;�+&Ludn��͡ټ��"�E���\�R#s��N)��v�����&Y@�H=�pY��faZ;2p5dS���j�9*��r֙��b���#S��W�Or��>����K;uk]�,��^�k��S��K�.��f�J�-��M,��CS���6��v٤�y�һQn��ug�u�������:'�6�<�\�O��b�Djܨ�)�_��GX�p/bYq�����?>��	O���=es��)����꒹�����j��_0�lK8hV�F��{��븑e�Ƃ�\v8�rNw5rb�Us�_X���:uK�j_(j�]M�*pn���ͪE�+�m����K��+&<���a@���i��`6��DA�&Y���Zߕ<T��:17� w���x��7�X-��6��,36�$�LL��4�0Ô�ߡ���1��8���p.�����'�6�ԥS�L��p��$m��
�,l��pbҟ��'F�?5��p2�v�_��C�C�ʜ�D�˄s�s�r�=�r��l:
�b�Ҿ#K�ГL~@!=y�� ���Ԣ�rb�ɣԩ�ù�bĄ'�zކ���M2�;�#����25�v3�>���|T��$�#GLĺ��k�^����0�'���o��S�[S1d��˛L�Y'D��%�_�0���@�� <,��L:��Ԧ��c^�S���|�epז7�u=��i�Ĉ��9�M��e�_�QFF�J�f�gq�Y+0b�H&Y��e�	5lVM��,��j��T�Ư}8�ɸ�M�k�f3��&'k<u�)�/�u��pY,�������|�{�������XV\?��s�ˉ����ȹ3����A�V&�.�<���S@�E�&<U��;*�2����l٘�wr�͍1T�a���ߪ��վP�d51u�Z�4'Fĺ���|Y�l̨��h.8��aN��f��+0gW���!f A�7�n�qCf�ސ�o�WG̅��
g�<�0ج�31u��Ü[n��'���1��8�H�\�=6m�#��#�ҩI�?�-�A��
�d�ܗ�YǕ��L�|��-��s׭�;6��7#��n�"h��e�nr��9X-�j|ҳ��Gȣ�)Ɵ�wiz��W�Ʈ�-WSe_,fVjy�Y91��Q����\z1b|=�<�޺�q�L}�V��1#�L-h���L��K��-79�E���u��r̀!��nV|8�I�4Ј�-u6`2d.����s��)��v�����&Y@VH=�䏇��?�Hk�q��j]�S�����ff�r�`�-1b���wN�a��^W5��([�+��U�K�V`�,��M�mdw�ꡩu�Es�W��aJ1�uk��>׽�q-'���D�Ӊ����pw��pY,KJ��~B��|�ٻ�B8��&bYq}ـy�X.'BX�̌�ې1S\�� Dne���Lﯚ��S@3K5<U��;*�2��R!Rٲ1s����ˉq�ͱyN�>9]�����r$��Q��͉���vh��밍5b~3hĬ����TP^"n���W`ήdݢ����d?+ݔ�9oH���#��CS��{�]lfb��sn���mD��c��qT=[�\�m�#��#�ҩI�_�&|RS�w_�u\i81���9��8w�z-Օw��7#Fx`��h��e9�9X��S���~�w�y6��5�#K�ГL�zh6�L��Zv�[�VjрY91��Q����\z1b|=�<�zPK��_�j�3r�Բ��M�(n��ȼ�m��Y.r�D��|^A`Ȭ�����'�����!S����%SdV�	��@	B�'L������ s�?���L �M�!4�u�O=7d��yp2b�,D�h�7�m?����9�����;G�4bܤp3u��x?T��0@��F���,�M@�u�#��n��pT�-�����:��R���l1�e�����p�N��������̷v��͡΁���W��M+I���b\W8��1�8\���z�T����Tolt_Ψ���~(W#�]\K�Lx�/���X�C|u���Yã��'�"���_!`^�T̠��Nc4�)�j�QS�~E��'��le�<�:��R�H�:6�C�^�0�QS{i�97���0��}�Z�ln�"M��y���&S�:r�3a*�f}���p�r��-B�z�9f���c&i�FќsK3���g�%�/F��8�WN�������uYh���F�Y�6&&L�#�L����i��I'D��%�_�0��Q?�p��p�Q����s�զ9�\���ޑb�W��=y�$y/�:���rH����Z��qs@æ��:3j���9�߮���f�@�5j2r_7�X�p����XW����~�E.綇'�B�f=�,G��*��W��<5w"<uۭ�&��9u̘I����ҍ�Yjdb�;ͯ�R�#� y%�����Q��o�6�-��=̾���f�nz�`c�M�z����3�E,+��V��M�+2�In戗s8�T�s��8�uQX~�0�\*'��4������~E��'��le�<�:��R�ȝ��r�̢rsպn�F�J�����n��"�����
��efo�Մ)��r�ٓC�~u���	S������|�qҷuw��9�l\��d��e��46fA��Kt_�1���Yc0|�"�e���+wH_VrĄ'}��i�6�4�:)��v�����&Y@�a�0\n)��22�b�ٸ�jӲ?�\��w�-Z f&�.D,y/�:���rHP)Z�;�|ո9�a��^�͚��ˊ��5u���jĨQ�"w�����u����)6b������I�*�q��b�\�o��l��;���V~p��:f�$��RF��`Ƞ9��aϾK]NA��J�1����&����f��>��:8\��������6q��>1��q���8��B��uEC&<��s=�N5f7�n��	�D]���+�+��	%&M���8>կ�z��$�������^Ǖ^*)ro�zl�΋��U�-�+�LLݢX�sc��a��e�6}(gfo��	O��E���fO�b�Ց�΋�L����.3+��=Nb)B�z�9f޴�b�$-[��ؕF��L#���b��#&�p8k息Sĺl�=������	O�(|'�*mfi�)tR�	��@	B�'L���iF� ���9(�y"3p��eW�����¼�d�,�@�<�R���CfAg��v�A_$G�3g�6�e%ݜ����]��ݜU]w6+m&Z��ZuL-�OŔC��_��p��[�j��,���ȱ��Y�jn��:2b�W�M��e�lج5��8LuO��dVbE�IX��A`ݖ��.���2g�K�L�m���r;6�&Ywϯ��~*m��3f�����s�=ӗu-;Uݬ��}�I
i���YB-"��[��5X�H�ϙHu`��%B����QO��A�6��ܜ�<��I��n��� �Y��&ƺu ��~۩��'{ҋ��l"�e�7��'e��b�n<��d��ṥ��t[���m#�Mߣ�-�sjY��R2�t?B��	�}1��d�M?�4j���&���n]�#v�WDLt�)��V*H�<a�d���9��a���[�U^�U�Mr�������b��ߥ^�d�
�˔��dc&A�0����ug#fD�S�΍m�T4��6D�B�nk�f��dM_�8�6/�F�M�<�:�pb�ֈ��8�<��Y��c��	S����fE�IX�n�dܘY�k�L�	3L_�d�n�Ews�j�$�_>+�lX�� ���[�M����u�-��-�s�M-#�.nV��X.�l�Ѭ`5-"��@)&*g"Ձ�J�ubR��o`b�2.��Eʩ��r��9������:&�D�˲�A�����A�����鱂օL
����JPn��]�mĸ��{������"��L����M.���l2���C�8`�D�?s����_1х��"PXA� ��I��>�h@^�lԠYzpqrN��$��lo�~ f&������dxd %��x�!w8��f5b֝���JL�:WϽ#�a�Ys5�&l�uf6/�IR4e���g�����x<P��:�9�o�0�=�F@5+
�Mª(uËuscfmU��h��5L_�d�n{6{��"S�&Yw�.:��r*�޼���:�IZ'g��fA���yݖQ
'�C���Q�b�9},�"Ձ�J�ubr��i4�F��
�w�n�t<�Ą���.�f�D��Ə ���A�����鲂օL\[f�t����m#�M���-�s�q��� *�����b�'ӫQ�G�8`�D�?׭�	`憯����S�	���3T v�����9>��É�80�n�.ƆVv�@] ��[�ˢ�
� T��VhZ�����7'���y�26�|�gr���ů�u�9�l��ba5f]�,���,�1Q�
�1fBΠS��Y9��M��9N�y�`�$H���&٬�A�FM�nѨa�����D"u`�l���4���s��٨��f�tݭ�7�
�O����p?�ueӲ-+���,O6pu�~�7��ycԺl�][BdĠY��O��b9�s�Y�ɰi��13Ú��5�������^�����Y�]#7�)[�`ƛe}:�I��n�8_�6.&�u5�pg�]��4zȬ�±P^g0l�eKu-�u�Af=뷪'�2?�c�"s��Y�wӜ2s���;VJM��V�&.ʛ,�Lĺ��Y�r���'<����yٍ�xu�W�����}C�^��Y�שӯ�ջ�K�L��b��Ծ�B�1������@P���۽�LM.f��i���d�.�ż.^M.g�k%gunzR����H�����j�M.{61e��J���2�zN$7�5aI�fю=f�ܒ�ӱ�� �uIu�ԝ��uY��O��(u��z.(;�$�Z��H�] S�lx7�##&��l�j����.~d��&Ò~؆�0�?l��+M!d�>��x]�fH�i5�$�n^����<��)�+��v�����&Y@̼���_�u[[5O��	���$��М����]Vk��+~�ܬ@9d�0n��\��R��l|9%ꖥ�W�M��-1��,?6h�uK��mU�����ں����a��YH٬����x8w�l΀d�z��M?=�D�+���˓�4�z�~�?(ms<W�(�,���&YwX^VlVo;2n*�V�z/�u2�&<e���fY��$\�R7�����3x��l����xP�������:��8��<��_�df���k��͈�8n�Ȩٓ�<7�9����t���a��x�n�3�2�6if#`��Nx�/��>e7~����a6ib���1s+Vw=V�M�_70�hଐ$��#�0rn��Zv#7uNǸ�fՏ5h���T8�bY����ug�UZ�&�s��ͯ$�ͼdOñ���HXGd�̧�X���c�209rN�����^�n�a��-�>lN�c�MR�(u'�³�C��I��]���K2�an#��
k�}sd��Q��9�"�e�@5p�8���7s����p���W0�$B����w��uUk��!�'9[%�N��]�������"Pہ�
�/O�d1��>����V���A�6�I�ӡ����cf-'8.�Y�rȌ`�D��ͥ����Y��$���p�f�]ɪyԁ��l���r�M�nu���f�Y���[{or�Q�u�A�B�f]�u8\��ù�5`�S��uG�M?=�D�+��ۛVV�!]x�o��z`�s<W�(��DM������8�ɸ�h[A���Ɍ���ƛe��4L��^7�9&�jR���q�Ñc�����<�2�J��&{������o�o��.!1)�/�e#�f���iN��l�L�!8NX���v�Ř�X�Y}�l�ay��	O����W�����Iʾ��=�z��N�n`L�,O2I*�Y1`�,�SI4Fn�l[�p�ĸ�fՏ5h�����ZH��I�]���.^M.gi��4��|��6�p��]�T[�βgS��x+��p��e��Y%9'������^pP0�[R}:6؜^r^�T'J�	��l��|��F��d�sA���j	����
+�]�##&��ɽul�D�ˆ�1�θ g0��篛s�Z�տ�_ס�
F�DȺ����͖�Z��I>��*��(ub�_�u�0`���8!�(A� ��I�UY�>����V���"^�f��&9O��=��d��y�ͭ 3���e�f;3���3k9/]5��̷�ud̬ہx1�q��:0қ�f�ۋ	dl��Y2wi��a��(���*�*8с���FΠ�v��|;"�I�av�$@"Zݪ��9���f��E�;�_��ɠ�C&ƿ5��»xwո����s0?��-h�q8���\7q7˟�͍QO�M�c�깑���i�3 ~(��S&�н��P1���-8b�R2'uZ�է:��i��4Cʒ�����ь�Bm4�z7:I�(e++��Z��DN�퍬@7���M_5�6�:k�Tr]�4�	�LR|]���!��c�ݸ�0�_�6��ck1���9Ѓ1�*1j��\�lNݤO�e�/搾t٬�3�ԇ����*K��6q�]��1qƪ�g`ਁ��p"�e���J�a���J�U�s��:(��v�����&Y@�<Bj���C.u3p�&3lj�A�֓ɸY(����py��A�|mW�Ѕ&�Bĺ%����͝��E�u_�d���cڍ�p ������KW6��?5\����AA��p�_�% �������$fk4�GL
T��6��h.�SÌ��Q��U?G��� ���9�,���+�֘� 2����������[=1����FNĺ���o�7���	O�Y�>g�2��u]�'t�,�O�c��[4C���&�w������ r��Q�V�в�l��&_��n�_8��������~'3EH�u��p>6�ca:��#��n��[��W��F�Lx����� �7I����_�!���Rb�$S�Yo1{��+�� 8j^'b]�3���$6aJ��dZ9��L��"N�@mJ*H�<a���#�fu�n���R}8g�6�� ����ɜ@�Lh2��L,�.�:����&A�huK`�6���A������.�=6Ǵ1� �u?6W��]R���u�.K���� �L8ҿneb�2�����,1)PE�[�M,$p��f�$��P�P��9
���:�~�OF8�nA�9}�7Nf�0~~4�22c|t ��4f��9�
�wW���Ą'�R��ʯDs�W���at��Љ�(�>�7y�G3�,�Ѡ���}��čNR9J��Z�7�\�H}8n��Ob��	@�Jn��w�1S�_W�;d���ps�0��˄��[��W��D�Lx�Ĩi^�9��q��)�l�7�,�+%�L2��%���[wM���j6 f8�Mĺ,�����+��Mx�G�+�VAν3S蠈"Pہ�
�/O�d�o}��r�`�/�'�s��aS�r+���G�l bf����Zz�|�5 ��V��K������t#n���	�:1fȌ��ҤeQ|�+�20n��:.��-<~�������t�rԤT��_Ժ �5\�lr��ɟu���'��E�O4�"�'ZYTq��������_�⏘崎��Ϻ�����'Z]D�D�-"��E7�_a��Ο(���?f܄��,G5j�q�- kff�/5�d���:��"G����UK�ͦ�$�D�Z������w���g)�Y�6�NL����µA1hjz3�W26ɲ�vٻ�s{��v�f6��j�5j��n�ذYH��J�I����J,�E�ݢ�L�(����.p��e�f�7�z�I��k��YS�e����Xx�xE�j-�5]�����[�5ـ��-�h�ɗ�ٷ(�4�lЬ��h&�ݷ������]���n�� '���J\��N�к-�w//��d��^r��+�l�D�&F��p�u���uKzhr̰��C���g%�+ܬ�-Psl,s1I��L�����,�Y���3S�G�;qܘ13���տ�gf`D��z]�CL��33����N��k���;������.��C�&���Lf	���,���sr,26��Kz�﫯F�he95�UX���7'4�bU�:7b��ΙC���j��u��G�I�F�r:3�D��>��l�:�aS�߂�h����l'É�,�T0�B���Š��q����Y�mjo-1�|�����y51��Rw-�lb�DΚ�9�p��ʦ���$]_��$�¼v+�,|�R��"Pہ�
�/O�d1s������®fPa��s�Mm��Y��)n�,�fz�pQsx{�����0�\ĺ�Uj΄uW�a�uh�+6d �}x�.��bws��X'��a�,\���7c̸�161e�:���.s��.@kFM��֍0h��)�G�[wb)m��2:�nS�����52���-4l�l0� S7-�f
�쳚�Xx�xE��m|Y��ڼ[M�m�#fe2��*mlQ�4���4�|��07eK���u�uj~���3GM�e�����g8�C붜��nq
tm�!��1��>V�9\o�M�Zn��:ɹ̵nIM������D\�.0Un1��cc��IZw��~2���,m}���}fJ��uh�\13�|9�!S�[zfFĘ����v�Sa��̌ ��L&I�vo��=8p��+�B�ѻ\�,_#8f���\W9���X�`6��M2�a����j��e0s�-���L��FY�Jb�Q�F̂t��93b�t��Ss�{Eo8��.�,����u��ͭé�dؔ��`,Z�4/�M�Q��o����ɢYO5�g&��Mn~�+�x��.[V{+h��9��T��l�\�ͫ��n��#h#[4�$�d=��ީxЇS]?���~61����2�,|�R��"Pہ�
�/O�d1s�����9�*��Y2ˑMm��3��P�q�0���f���x�b. 6f�s���W�9�]M
s�f#3 q��T��-����!>b��R���gf6(MMof�Ս�I��q������NM���s�v�5�&Lu�v�+� ��u��N�A��RJ��:9�6ww�F�_�e��͑&%�-[�6�fQLa�}V��a�LR������!Q���[�5!#F��,�)!F�M�-�%�M-#��*�i9	����OL[��]���ew�Iq��U]w2�g8�C붜���8tS'fȰ�d̀���f�ہq�!0�`��\�Z���&w��d��>W{ۅ��-f�vl,s1I��mO��
Nx��'���g���^��uuc�/'9d�n��Z�z��y��
�]gf��_e2IB�l��܃�ʿr+t1�h�$Y~ޯ�j-�u�S��
9'�5l����0~O��e95�����2�e�*�	G����9���1t��k��,\���0����m4b"�e*/�dМ������E���9��{�4L�\z5�g&��Ǎ/��s�uٲ�[A�G�)��Ge��o^Mi��A�z��0��ܧ�ANu}AY3�~6I��<�&���v+�,|�R��"Pہ�
�/O�d�_}��� ��
��Y�ˉMm��3�"��7��^�z�،��;l6���fs��Қq9�\��2�Rw�O�Å6ޣ��.���!t�a4�u�$s��QQ�տ�d���$�Lx�Zw0+^�"�E4*��0j�� !c@&�1�9讖4n.݈y��-�M�$^����R�_���Φ��.�Cy�w/��!s[�f
�M�����e,�ӳyj6��̽�@?un.����r##gꖓ�-�L�s&]_PW��ը!����]L8�n=��.�ř��
��Ǹ��+w���6ɺ����Y�Ņ�2�_L+�
V����2Y�"�ʭ�8���I�6�h646c�M�����[�E�(b��EZؗո�u�����f&z�:8�=���M]��.
�B�.�nb�.	abB��,�_�0��u]3ŀP��(��-'2��j�Y�*⢽#l���L�);Ѱ��JʩD��Y��J��dj9Â��W/w2l�1��������?�e!�L!6�e�݉�����Q�(՜Fn*���8��p�!�dz2��0��i���A��-���q�Ǧ1�V�b��-�J�����Ͳ|�V���22WRM��6���py�)�G��o��N'D�B� f6���K2��MJ�p@Mĺ�Y�e&�y�2a%��؀	+A^��%��qx	�U/A��愗 �;E�J��-��%��&��F��d�l��"O��qa��`�6+hTӂ7s_��߫�͟����n�X9E�-�a� #f%�$�N�,��;�n�z��!��;�����%c��N�5Y���Mf��-ܛ^��aq�܂sۇnbꖯ�1�̂�����&�}-2�_�f���M=��ne���e�����]�%�4k��U���:�6�1Yw)[f1J�����s/)��.�[t��i���?_��	����q�ȴun.�ɦF��c�3�4����D\��^������;k��l!2SquD��E�N+��͠��Y_8`Z=8�r���Ir́�VmrY��u�
Z��z7x	|5jj�.�+`���dݢ��+w��1S�[ ��9)�L2=�{|_l5+���/���L
Ѝ��[�q#���F�Y#0r��I>D�I�����ڿ�D�6�tg�Ѷ�.��,�Y,ndΝ8��9��I]w.d`6��@�����[N�ͦ$��ɴ�h���]6˨
m�ݰ��i�&&���so/����vHVs�_�$��}��j^������s,�TLك����b7�WiY��Y[41�-g�f	�9�n-�.���$d?'����ɩeg��&��jVК�YBi15��Z��t]cd>�ڧ�=n>��	�ce��ph���i6S����_hpb86:5�A	B�'L���!3-?�h?�!�N�E�}fS��&���)f9�fp�/�h�\�{�b�̨y	�a`�׹R=���X�q�Ĉyɦ�H8��hĨ1�&��U7}/ͽ&c&ZY�I�b�^b����XVR�p����>h�T�X�͞D���e�f٭��ah�-v6k�F+�M&�Խ`Sp���J��҂��Њ�IN��QF�!L�;����m�����Y��y�t�e(�X�faZ�봒���n��K�L���	8C��4C�q2Pu�}���ej�ݳG����L����c����0�X�}Ǐ(2�\0՟�fs��d���v��?Vk��y�\X73I(6h��ɈY��_p�ӲY�d� �<
�N�%$��n^��j�ؼ2phb2D�p8�#31G(�	K����Ir`џC��N�A�]�Rr�܆��j��7��W�.����Yv�fsd�	S�3�H��+/���̅�ҵ ��Ã��gy�j�N9#������ -���M����S��?4����ě;��"9��͙��k�(���H�.�q�#�e�nؼh���	S�Y�Kek6k�:l
)��v�����&Y@�4M�᲼�~aAs�4������$gy�A��d1dN����dL<��@�jְ�&z�j�y�u?D�IAw�/��<ِiF¹��F�3[$��'9��[pȘ�VV|:�q�H������>��̢:�4�\ϥ��45dRV�lY�?�47h��������o �պ/<f�l
��v��wioÂHFL2�1�����,ܵn�W0����R�������n�틾|N:5w!ER�:6���>����j�܃-W~��I��f��j�!�hX���U��f����gޔ�����hU�'6�D2f�o�XV�"���.�.[k6�n�O阺5Z�#�� �Z�^7��Fh�$	u��Y2b���a�ͲY�d�������>L�A���7p��"�G����|�"��e7a �9I,�53d_��4���+%�mH�}a,��zSᨉX��-��}�2\W8�I��U>���R�`�B��$�߄����m�U+w��-���$1h�6I��(���ΝO&^rh��%��7ܜYk�會��1�lb�_�movĺ��1sm�ey�1��8����-<k�:l
)��v�����&Y@N�z��r̡1s,��f��MmZq4[�r6�,�Ylf|�o��+���I�>D�^o4r��S�fӫ���<9�n���Y�������4�w�9�j��=<��v�f�QS��'*���9[�l/�>7r2����r���9p"�e�Vq�f�,L/$����Ss��h�"��/��^H4`�T��Rg��ί��e'�ɐin_r�LӲ^����j�9��i�mnc`?��M��6�ۻZw�����F�̷�S���r� �
����
0����u9���F�z
7��#3�.����0խ��\��[��Lҿu�Ko�beW4��-�|��Ij����
0?���U�߲�}Y�As��ہ8�p����9>�D�K�|!����b+z�M�qs�k��9b6y�0&I��_�Cٕ��~\8ԭ�"�0թ�3l�+��;J�1n�r6���M�_*Һ5tu�z���Ӂ;�ۡiMW��p#'b]
���y�~+�&L�"�˸5��[�[i�m܉:1�t1��A��,���}4��4-��;h�)֝Dg.�蚋��Tl�B�RO-�`G&�^k����#SY�և�3b����\4뻲�G&ZY��hRs.mx}Մ'���K���X9Dnz-�8�"�mz���lF�1 �����0�1����6XZ?7�4h�ގ�hpcfy=�";���e���*]�Ep��'uN���h���qS���"Pہ�
�/O�dAs�� �e-jF��y&o��6�#s�e۬03��ɜ<�Vn*�Ӛ�9Ö��dS�N�5�Q2�Vi=Nw6`�d2v�
B�ΛX|�Y2�v�٨�-�C8��p}�Ԭ�9��n,28�_��u�77��C��	S�#�p����:���x.4nиI�7��,Z8^p*�/�k~��i���n�͸Q3� S���O�2?��A���nZ��w|w�\�e����hi���Zǻ�u�q��^��ˉ�;&��S�.�}ll��,o8n�֕������/U׍���ū#&Lub���9�&#9b���;MO��@:u�|�m�8i�O�W��b�$�w�w�c����s��N��i��>�D�K�\�1���Vl�!�³LȐ��[u��#ƌ�C�01�ZK�Pve+�W�-r��'6h�T��k�� ����Q��l��*���:q��Ѡ��d��l=֊������/��s7�ȉX���f����fЄ'��,
0�~j�]�~���Aq�;Q��	ż���`^���дp�CbF35�Dg.����Tl���S�9ؑ��ԩ������TV��ao3�&Iثff�Vv��D+�~-�x.mx}Մ%��q��yA�b�T#f-�A�R�:2��f3�(uf�.h܌ cX�H��XZ?7�4h�9������Yd�w��l�������Q8��3��{��)�T�	��@	B�'L����}���5#��<��AS�N�����g�6+��7s��ɳ>�}E�rZs7gز�����9��А)0���X���S2N���&V _�j.�B�p�I�z�ad��P^˖�Z �TN
�SǦņ�����X�}�s�0��z]�0��C�ulਹ��u0Kw�,\hܠq�L/gѝ� ����5�Z���X���q��͋�Ʈ�&�,�41�/߂z��]wWr�nvuR������i��w����,������Vs%7����uٿ���z�Y�p�D���Őqs[VLͥ�qu�xuĄ�n+w��*5)����.=9{����@��u]ݓM�q��P� s�ŀ��4���X����Vos�'N��t�|��X�`��cͽ�؊��� 2�tqv��#ƌ�C�0IR��!�Pve+�Wlsb�,�OlЄ�N�!��\7I��ԙ�܁U����M�09����e�VlO�o�Z��s`X{9�Z+�Ɲ��hM�үߢ]�8�Z�w�J3��$��b^w�
�Y���>�av�6y�����p�ሉ�Tl���S�9ؑ����	pΑ��^���f�]Ma3S���G&ZY�k��si��U����^��t�*VNI5b�R4q*E�[��f��Q��]иA���=_�����)�Y#0���c��A���,�G���x�+�I�fn8��{��Y�qBj;P�PA��	�, l�?�pY�C����:s�AS�N����U۬3��\�,�E8�l�M���%g7'���Ь�F��� 4�R'�tXG8G��J�mj)���r̠�#&T�̘YԜsjR2F�,RY�˳<��0��<S�h�<�"j��5@���(OԺH�D�,(�c����+Ϻ/j4�'Z]Tm�7�'b]4y�Y^y�� خ���w=���ļja����YDdB�n�шa�fO�H�E�/�NLX���9��l�y&��_p����3�f��	#^���
#��E�OT���'j]4q������ͷ�ğ��^��n��˟�u�ѿ���XQ܈���."��^��M����|�v�Z-3p؄��њ��xF���#�f�u3~�I���g��ll)��er�, nȬ��m�V����]�-��K�Z��s���u��<+ef�@����������Q��o�f��f!�S-Z�g�/������q�����I��.#Ǫ���)��4jB������T�-�-��1g�c�]���=��l����e9�_C81u���|k�TjF�KY����Y'6d�t��Y?8Ef0���[�b؄�n�~1����Z���rG@@P���
ݐ�0B����	#�G���]��Ąʧl��N�|���ʧ��	#�O�z/�0ByԺhP�.#�l3l���#�E��eѠ�����	#�wݚ�	#�O���F(o�lZL�<j]4(�XY�(NPnf9�1^(�2/�G���/[�a��] a���-��B��.2���m&�P�."�G���ȱJMX�<ZYD(�X�G8f�寻��
�S''�P>t�^(�Xʣ�E�;���jP����f6��׷ͫ��_{X�8|�����ٱ��q�20窘�
0�^8�����Yd�Vf�/)8jĴ_�k����7Se�6+af���y9u۞�����ț��2s@?�А�X�ӯ׸����0%_P���ň�S�/�cwA��1���r��36����I~�cҫY(Vb�.�p�Ժ��V�� #�M2������YM6Ev7˂���:�T����Mf֧���dp�ﭙ�nōas���w��Z�;��8Y�|���A�X_���Z��C��Lx��M�8q���Ņ}���L��@��!�vv��M���!!��ԭ�f���/�M��(u��L_��QL��Y�nu�,�V�̦�\j17�M�6u@�s=ؐA�.�}��y�#���K�6�Sf�|�x�f$�ɺ(`�~r�L�-i]��e�f��n�,�A��%�N��:�Cיa��Q�⊁�Km�ù�]v_�i��$���[s�x"6M����ù������h�d�`��e���OՕp�M����\��5wy�(�ް�l����)u�h�u{81��Y5?.22��R�	��@	B�'L���9�� ���73�d�/�۠f��&6g��C��ݴ�f\����9q\^]0�ăh&���<�"�f��A�&Le���g]��
)p&����,M���̉��:�_��o??o�i�"ۚ9?W����t=S3N�N�5皛���u9�23�Cfq�	S��=���������F��Ƹf�����]�Zǆ�I~Ó��,\h�LӦ�-`+�*n�zl�/���ա�M��Ͳ �D�!���$���� r���m��[31��b�3n��w�@���L��Cf�C�X_��z�恏�0%w3Dw30],Cs7��K�Ab���:��d*��Gܐ0CJĺU��ѳ�n��G�[�����11��1`�l�f��jfN�K-�s�-2K�\6d�D��|�ʬ��8�Ò�D4��S�����e�#�uH�E����f�hI�"��38dv�]�� �>�kq���:t���̨6�1��+r̋�e�e�jN�H�����&�z-�M������p����kA�Z�9e�Ew��0%_�r�6k��Z�5wy�(��㺯��)u�h�u{81�:x\w8���j)��v�����&Y@̜s}�Წ��1�L���j��ibs��94n�MKhf���\l⹼�`�є�뺱���J,9h܄���5^���)p&�q	��_�=��\��kw����Me��%�)3�}U�Tp�����k�&���N�s��ЈLĺ�� �n�Ą)�z�����{�u���F��Ƹ�f͖�񵻶�nSh&��Ir���M�[�δ����L�߸��:�ɦ��fY�Y�p��t2ɺM�9�"��;�Ԝ�]�f��=׉�h̸����ٺ0S��Of�C�X_������O�{�]�s�-Cs���LA�uj�m� q;�N�a����nU6s���C����Q���90+FL�k�FG��_n����5s�������3`�_�s>b]J��Z����ux�o��B|N��:2�1nF�됬�6�'�8ђ�E��g�ϕ^��m"���xʸY�u�:3�"3��Y\1p����H��]v_�i��$���Exz\hkф^�e��UR��$�N�M�d�`�����0��J8\��%=X�S��j䨹�E1`Df��;9o�#��ݣuX����`�By��\d6d����"Pہ�
�/O�dYǋ6.�z5�,����o��qv�؜�f�w��y����β1s8�(�%0�yo�KZN�y��9�$,V6���}+Ef���Ey����^eB榯�sg���D~��y\��k��tY�TL��1�A.�*��լ9�i��ŝ�t.�y�G�uKxs+xMS�N�&̨s��n���j_37a��);|�l4\��̦�⦷cS�ol��,�;��ع�er��
Y�;�FMRH7��~a��W��\�]1h�$�~������K��ͬUR�Huwm���Ш!�_|ݖ������T/R� ��(�:ddN8��u.�i���I~
/�1�o��~b�tSy��,�jNT51��R�Y9OA&Le{�������5p���I:ݣ��.L%��:���j�pj�Kha=��T��qY=�?2C(00E�������C�Q�I/	��~�`s���2�I�_�ϭfu�&��Z�\akgfb��gg�;D�Mĺ�~�ù/�ڹ���E��|%C�Lf���n��^�:7�
_��5���Rw@*�5rb�1f̠ن����8_)7U7b�w�҂���t8���R�L������/�U��X�cq]�y��Ksu=����:s�{�_'F���V�)�ИDn�İ~����o��Zw�[I1`�e���Hu뷂n��$'Fx�l��2cs�q�un���eh&�l��/h�D+K�j����J��莞����1s�D����FӺ�Q�L���Ρ	M�u��=9�ԌgaQ��^�+��jb�t.���V+%��'f�g���ĸo���[�r�n�-N2��&�bg3p}"ép|��96�l��/���!��AS��.�>Jn���m��Zv�:ܸ18Q���'�:��q=J�����jVD���,�b��o�e�&F��\�`r�D�Ks{�,y8r2�DO/�$Z�_7n�~ٸ�i7�AȳMғn)Ǡ5
�N�uY)6ת���"Pہ�
�/O�dQ�����'*3j̰Y��S�aMm:l��jo�ͣ�b���tq6q��Tj�����ĐS4]|��2�gClnD�����ٍ�!s�&��s�,��nМ�k�5Y��;ٮ���k��=C7}�ǔ�B�9����j�i��	1uw��=�F�Ժ%����4i�g)��x�W����F��u���8uk���`l�D,S��\a8+���W�K��uL��n/�nn���&3p�n(���p���{�s�٨I�����
�����upV���l�&x׭���p������lv	�YY3k�Z���v�WneՐ��/�n���v,Z81�E�S����� '�ߡ�z�9��T�G��O�&��'?�O�`י1��.l�SM���r�<�0�]x��F��/0����2W#&��s`͇�`J�u(YJ`��qj���2g}�u�3h\V�����[���U�����zˉ�6�����Y}45����fN�I�_�3H�v+M���ܳga6c݉x ecf�!�&b]��u~ 4�1�H?�r�,��3��Wc�BL�^�:7r�\5�k81 ��0T�j�Ĥ_bK��HFL[w����M�{ݪ޺�Zd�Tt��>8Qj��n]�}��j�M�cq]�y���w���p�aS���]o0g�fb������5�S�?f�[41����[&g`�;ȭ�0۲���(u뷂n��-'��#��]B����s3�<�_防�G΄"s͢�%Hef���ڨ�莞�R]6K�f��>���hZ5j���j��Є�ʺ/�{r���¢ҍ5s`?bդX���9f��T�.��@�&�}7���-{1�[�-�5X��x�1��������Aαaf�aJ�n��ŏ��K����t0�4|�\��t�#���Vzy,�8��Rg|8	ׁL��Q��ܷUV�"b�Ĥ�`�1q6-|[.c41�]���p �Mĺ1dεeGN���՜DK���­��츽i7�A����'�B��(�:�e�؜S�mE���� T�~y�$��&�0�S_�B�Zǧ����t �������F3�̆�,�M�q4�j:�r7���ɚ��p�����kv��d�\�ɺ���e�PB�As��;Ԥ��nSj������~m��M�1e��
vs�-l-���_�"'%��m��=��[���"b��$_��^+f5��/dpκ�H֙9RЬ�5s�,�u(>4�.�IN���f0e����?d�~7)_G�EY텛L%�V���y6jR!Mݙr�Mj��
9�.������.�9 �1Sӫ9V����V�j���&��RE��LҿuG=�mo���IՋX�f}���N�+��s.��P�����L��W�|?1�]g����-N5	��w0+1�_��"�21�P�ʮ����&�,g7�\����3s��)ɯ֡D΄K95u�~��!s�W [8��e����ܗuY����\�@��ʉ#�yR3����_8�ܬcv��$�/�3H�aa���ܳ�1� 9�m�/L˙Mĺz&�:�pĄ'��반ќ�dȘɬ��-b��E�[>d.���5�$�F�; �o�"MZ'�V�1s����n��n��	oiߺ�Zd�Tt��>8Qj��7���6|9]�kr,n|�'�_�sf��Y�l
X��뽑����Bff�+s��T���A��M�S�[&g`�;ȭ��� ��u뷂n��-'�����6�7]�f�yX��1$ۤ�	E�E+K�ʌ���fARS�=5�{�,��	����n�i]ԨI&?m�,�C�
(뾌���f<�J7֌�A51Xz����J���]����AL��K��-a9l�T����M<t���N���c��&�/�+u?�jW,�6b���P�����8Rk١k�ٸqc&p���N�u �z�:7�m�լ�61�#XvL�Mߖ�ML����۞,n"�e�bݖ9l����x�uS�V�Pv�޴�� D̊Oғn!�Akz���RlΩ�"N�@mJ*H�<a�d��ս����f����Ԧ��t�7���Q��C�0.p���WyZ݂sʬ�j��  �ԁ��̼�Ȩ"ù�g]�,��ܮCs�oҺ�)��4h��Y~n��^�����.q�gҢ�,�*8���;B�G++>-�e���
�
Sꥻ0�a��T��	'���M&�������9y7��Y ]GH��R����$e4D���ЩY�ǔ��1|�l��Ϸr`Ȭ!5n�d��.��}w-���<?Ը�d\��xٟ�r�����}Y�R�fi��uݼ�$'��0px@s�[n2k��\��,_3ɺu9ho����Vm����`�X�y��cd�FG�ssO��BC��{I,�l�1�)��/�(a#f�.F��xt5�U��6�nf���3�qCm9`�#����P��{ �4Ȅ)�0f.�E���4dnn�8؃��C������ɬ��ڠ��&�l�jK�$�����c��ĸ����:V�+�F��a��z0SGM���Ks��sĀ�pi]��15���!{�O�����վ��Z�����b�1B[��t����u�n��=���܄'��Ɍ��vV�n�!��H������e�`������n�-���13��=�Ay��Zw~/1jnS��<뺭�7n*ˏ��؈�#4FxQ5�Va9�j��]6I���4�'C��Q�l�*��h����o�3|ٮњ.���Ѳ%s
۵nY<ﲕ3���˷���������Q�V�2_�N���hn�Z��x_��!>Yw/�纴j������Wn!Rgwm�D�ˬ&3�\�m7�&<��a����֭�57�y1ۑ)�)��v�����&Y@�z�}��
<��Y�E�d��6hj�j����v��<�J.ǭݸA�f�L��=0�ڗ/�y����_!j��:7W���i$�uj��9!v��/6�����dæ��a��Y]��@9X��?SEfi]��S5�ʲO��_�+-'L��0`n���{�>��!�L>=Ǿ�E�}���9j:B2}��scFf����\w�P�СY�K1�}4��� N�WΤCf٨q&�W��q�\�Hl����k[	q��9����RN2�6��}Y�R��p���+�ᔝj�b4���&�7����pf�u�r��(�M[�� �1`�X�y1K�L��Q��ܓ'�����}"�9Ĭ��꾜��Ͳ3�ujJ��U^U0�o3�ff��ʸ�����q=G��>B]�o0��%�ؐ	O�3�e��m�\�[����l�q��F�As���d��� �4r�Ĕ���t�$����̱uib\����[Ne��r�-��g�%1�ީ��k�E�4W�?G��9��e	���������ʧsL��}�6p������t���a��1��:b]N�5��t8`܄)=7f��Y4պ��!��H������e�`���"�]�����8�����R���Vs�ަ��o�9{vT8����ڙ9Bc���od�*,GS����ƨf�~⃁�!�̨s6mC�g6sl���;×��|7I�����L�B�5?,.[9L᩻|�����@�p?R��]�+�@�I�Յ�DEs��Ժ}aY�׺���W-j8�K�v
.�p��47'F�8��Mĺ,;�����̴�'�&�9ԜMh1+��
�����Z��"Pہ�
�/O�dA��>�pY����_��Af�o��6�������+5@�Lp2\N97n�� ���.�}�R2��6_����M�� �Ϻ�1�H�u/�sB�.�j�ax�]��,?7�a�~�,`wg��cU� `�)�j��1s]�l�&ZY��\:nNͺ�)��3�mAVwo�֛��d�ɏ�+�"�r�l��Q�b�G�;7F`d�)���Q�j�\�������m[
`�Ty�Lj0d�j܄��]�/�@h��l���y�Nf�TH8B�aM�91,����u+el�K�8|�f�,7��-71�;>3��L�n�?�o���i�� 8�X�y:2lIףԹ�'Oz��I�}ﭘQWLuͷf�,�L�d�Q��}8�
��mf��,?8C7q�5s���j�u)����R`C&L��Ϻޮs�!�̊l�pⰵ�o4G��NOfm�hԠ��&Yf�T�R6ɬ�&6sl]��WwSG���,V.�C�6qXZ_7�'Y�c����
^��H�w�b;3뫦�}�=d����~ν!j�������b�q�z�{礎X�����y�m��	O�!�=�6+��Zw�:���I��Ց1���l��1�ꮻ�M���c��׃�Rvs��u線�6%���C��7��G�*�Y;3Gh���n5�Va9�j��hR��_]8C|0p2d�uΦ�b��ѽï�i�3|ٮ��v��4�/35`
���aq��`
O��[���]3h��G�[��|�8I��z�OT47L�[��%�p�+��>v5�ѥU;�<����!Օ7���]$h"�e~��0k��iKz9j���@�YЄ�Bج�َ͋L�L'D��%�_�0�2����P/��_��Af�AS�V��Ȍ�n� f|�sY�X�M8m��������Zlݒ��pV�.�	���p�,hrγ��Y�rp8�����<�΁Ň�L�x�����B��z�ݬ��Je�Nݪ.����J��9n7�&���P7'��e�BƉ~�6���d�:6�����d��9��d�t��Bo��Z�j��L�$�Dr6�F�<�g�0�-��z�-S5���mk�Ҩ@�4lku���B�f�c��v@\�S�{������ڈ��oQ��.`�/�k&�x��!�� bY4Lق�L	0uk*FM	0u�vz�� Svwń� ���c&��L�0eh������\��`�6�^�#@�����#8�7f䄗 d��J�he	�^��\+^�FLX	0er�K��m,��:8a%���V����� ���`\^D�Gx	`L��̆��&�8ody՘+�ܻ�h�S�BN��DAS�n9+pSp�Y&Eө;��o"Si���[��Ʌ&Y�$ɘ�-�ʸ�����ĸI��$�|=�v�)|��[э��|��%	fY,Y0n
�_0WL΢$C&�.b���nsjج���oQ��ewH���������|A��u/��+��p�uW��q9��.��х�W�By�/;8G���b�����"�&���N�GX��^T��Vf�b25��|A�.8��
;)��֩Yu2��MÜ��Բ[�]71�vsҜ�:4r���2<RW�M�E��5��I�Un��16[-*61�ɜ�dN��2j]ʡ��H+�FO��a���@��,]1G`
D�rV�$saT��-7G'��P"՝�K{�&:�ԍ�r��A㟛.c�����uw�в�,�j�ur䐑s��fZ-2dĸ9_W�&ƀ䚲Y㕾j��[?�
i�Vy�% l@X_6r>-Í� ,Z4pn��Zw˗��A��1�^���]M�2E���� T�~y�$����cu��Y��y^x�l5Ѡ�Mk�L̜O��Xˇ^����T]��6)_^�F�O0'�1���v��`�Բ��0l
�6l��S��ʁ�Md*�8�X̩�&��:487d�f�rش��9벷�r¿e��7G��Z�f�Y Á'��<8<���[]���#g#�0,u��?��`9Iߢ�md�-K7p���|\_�6p��u/\�ہy�TSw��ك�D���-�C��W�B�&L��#�q���-���6�&�_י�˷�Z�)�]h+��hbX���8]��Z��
�3^�խ2l�n�
����{IV�_�@0�3l���Z7qpV�ܪV�qs�t��n殞��eԺ�C�����Cс�E���{����#PM��*�mא̅Q����,H+���J���[�
< ����(u���=1wM:���؜�`2��[s��,�j�u+��'feɀi�Ȑ��|]�71��a�m�j��[?�
iSK�Zd:�ۗʧe��$ \��GS�n�������c�ʊa�2��qBj;P�PA��	�, f�0\���6j��Ϛ�&4�i����S�	�l�
f&4��;6�����ym|Y�M�q��76
S�u�ġ�Zv5���d۰I�|ݭ��i"SYpo�,c1��T��-�=2�l�rش��9벷ŸI����wޘ�FM�[��}��Tx7ϫ��T���#��&<u��?�٬���oQ�����R�VNL�q}A��!�ֽp�nw蕓���U/9����X��;�͕�&L�lo�yPӋ��mn#nR��[��Z�)�]h+Cfu�İz4p��SU�\a'����a��as�uÆL�S�P��{1��̲��ͰY�nh��Y$�lTs.�Z���;�0cR/��z��Q�Rmvy���|�n��٢BS�=KG��&I�U[�bN@2F���i��`�B�Twr��otD���\�wM�nN��qi�4d����g�Ġs%feɀi�Ȑ��|]�71$��]�
�K��-��b���ޣYBˁL';9�pdb a!<y��抩u�\���R��1|a���qBj;P�PA��	�, 7�0\���&�u�,k�Zh�Ԧ5\�fN����ͪ�y��氵���q�A�o�t�sS\z�&����N�'�u��m�s��,��[���7F��{�f�h��mF�0�.�1}JƜBf��טu7����.�1�|�1����y��ã�
��ͭ!�eGL��bЬ50볻�fB�n#&2n�	NFF��Z=9��3h�U��r�E4�-�%Xw9k��/�ɺuc�^`�!��]��{�Y�ۉ�:1�����*݁q�u� sE��2��[�V��Y�h&b]6~e�}As�ш	Sz3Wq���N�oi�������	Sݥ[(��έ��n"2˲��6�\�-��MM��ْ��+wGb|s��)��d�&���i8�1��9�N��]Nĺ�c/:җW�/r���[��׼"y�.��}��u+g��`�lV�Z��̨������7�~9���[�`N�5V�Tm+�������.����}7bNfa��6��r�@�D��̦�\�1u`^�(�lLM����b�[�˼Č>���۬�钉�ncd�\��j7�2�V�hl��	S���B�rGY5^̘�F�A�#ԭ�����$��Rg�F�z\�1��հ9k਩[���́AM�V����f��h"������J+	�M��?��x�]�F�9���Y�lb8��C�ʭ�9�Ѩi0X�����������ÁS�^+4϶�u��L���7t�ќVG��'��J'D��%�_�0��Bש���:/t���j��6hj�W�f���k��bج 8G���u�i��w6���yq�)���F�V�{�C�n�W�f]n��h�Ss��ٲ\�͠	W��˸!5�ٚ�A�s����6u���М�lnv�[�x�m'&�m���U�+RE�����dR4M��9��,�c(b]��o��#��9���~��*9�ed��j�Tw��q�s+)�ub��5�#�?8�|.���0{P�F̕�#Iߖ�8��^'35���1��/�)�Q�.�6����b�R��Y�`�h���/K2�����]�~��f0b�u���J6̆�j3�Ҧ�b�nMV_̳_��9+̩��j����Z.h�1j��W�n�1��'��/���Z���Rs��],6�baz�N�𲖛Y]51֡ XbF����m��L�֭;��٨�a���uٿt�5YՄ+�}Y�y���aS��i0��i��u� sZ�����Q�̜�����c�/f��欁��"l��>351�{�wn��h"�����݌ W�0%�����J����sna5s��pj����[g5r*$/���Z����rs'�q8��ͣy�M���D���+ ��;O<9�T�8!�(A� ��I3W�0\���΋t�m�ڋi4������p��73��,G5k��+@L�����`q�ɮ�i�Ve}v��L�ԑ���p���߂��ٲ\�͠	S�F�,������ם��1�7 ��es�k�z��n;1)�%���m9����Q��K2	4M�6��euE��Ƴqs`s��aJ��6t �UX�@���&Lu�n�\�;���E�;��9V����`�|.���0{P�F̕�#1��瀼�GoM��h�,�{aJ��B[��aݶt�FNĺ��G!��>��_��o���]�~<2�^�:5'աd�l���ֱ13*m�*&����g��}7rV(�Sw��$U;�4h�1j��r��Xc8q?�9/^N���Z���}rb~��fQ������e-7��jb��nn��}��+�ًr0�����ffX�&b]�����i��	Sz2K�_�W6����s<�1T�P�Y2��?��I����)�����c����YGMEغ�}fj�H����f=�D,KI��J+	�M��������9@w9#¹���8%�\�uV#�B��h0X����6�5S��0��p�T�7���6��r��l4��f������59��R)��v�����&Y@�b� �0����f�W~4�����q7p�Q��N�G���;?��f6����-�T.9\���LF�!���;���hYɸIe{�u\ڋZ�-�����Wdݳ\/���뎦�~���e�f�p�:5��4��g&b]��H��l4jYNNf�X�nV����ۋ�̧����ES��7�:-2a2�����c8�Eky`:]S��0�
�P�&<�oj��9Ģ9a�c0����@j܄)�Bq��\q�f�7~��UN
뎭������$��P��f�d9�d�ep6{:�Y�e�/G0p.���w��Рٜ��Ƞ���TBs����6+�f]�IL
���'E����ur��9,�$db8��c��^y2�2}�7�3���?J�\Tf�daև�1�Rvro6���"�E��C��|`�px���p����e��0�-��Fs%�6�8�'���G�jʩu����&6��-����rr�����+��VvSp�$ӯ�UZ�e�f5aҪn��	�6s���3+L�W}Q�q���ɜ!s���5fԄ�n]�j�E�&Ʒu���ȸ,�K��S��R�	��@	B�'L���y�>�}G��N�m����ڴZ���Ŏ��g-�%6:�	m�Lp���r���6��D|��3!Rw��w5G#7l�u�t��0p�T>-�Mo $���e��fQn�q���ܹ�A6�XL�Ssq���u��L�:0�n)=���LԲ���w��+�fۊ�M�9\�+1nRП�۾���eB&F�n�D�Fp������+ef7��23OKf=��e&�^`Ĝ3w,L_4�@j܄'�;̬�D8���|�����'Luh���_���Q��/J]4$�Uj�L8�W8:��m�����nЈ	W4g���)hbdޘ47[L!�ځa�rj�u��d��)��:l�`�AS�䰑s0I��ph��Y�C�ʓ�X��/������0��ej�lrQZ���p�1�Rvr/b8h�,�rb|�PQX�'��d�7>G+;mB�
_n�	S0�Y�ݜK1@v���2#�֝�k$�p��
^��\Nn�T0�veɬ��M���L/�$#�h
�"
i��<�0�3����^#�0Efy�	S�,J7l.�̙%��85a�[ש�f�f�[����>*7�b�ȁ�C�8!�(A� ��I3O����:��Y�bR4hj�j���Y���³���
��q�͜	n�gg��ֺ����p�C�L��]��]��H��d��n�Z�l*���^�_���/;�.ʍ<Nq��{�er<�I�-9�뺬���uٷ��m�S���ͺ�YV�V\�a��p��hĸIA�ɲ_��mx�^^h�����b5��w��,�fR��p��˹���2��{ʕ<gN�p���]�L 5n|�&��k����hs#N��Ь��?�FMҿu�8V�Y�.�KD&:��m�����nЈ	W��<S7��P�&FH�6��f�)$Y;0��u]�"�^1l�a9,f�ԺM�Y~fF2I�,7���,�p�D�K�f�oz%�<h����������9��4B�ɽ��a�@ʉ�-B]Da���N�����he��M�Y���4a�CfABsԻ9��V���<��YM9���^#1��X�ج��\Nn�T0�ve�\���#'�~Uݜp�ES�]H��̀�	�������!'L��,(����'sf��9��,�j�T��S����&Ʒu��-�y7��ˁ�C�8!�(A� ��I3O��c�%tJm�Wv4�i�V�[���³�Z����s��nĴKf΄-��3Nvk��p.�]6!Rw��G�"Y��_,�n`*$,H�o�2�d}��[.|@1�ݵ3\���(&Yw6�9�n���X�}�_~KyCÿ0�_�r̘����D�c~Zbܤ �5^�QM�rt���9��֣�)F�Gͬ����l�MŠ�+n���rX5/;��}x�>���U<��	S�[�F�4jnnǛ��6LuӪ/|Aj�$��P�/cC�0^�p�A����巄ݠ�:4h�{���b	�.��̹T��5��f]��DJ�߼��3s����n9`ܘI��pj�гT�y5�R��9�,��NN���As�7�_8t!-��
�!7���N�/6�W���BZ�k���%x����Ͳ�s���4�0�--9#!��O�/ �`�컩p�����T��y~��������,Ě-�r�������	��ܬ 3�c�Vc�
g�]��5<(�)��a��n�Jf��E�,m3j�T��Su [�c��P��+�	�ɍ��S�8!�(A� ��I3/�0`��YB��6��.�ڴZ���9���f���j��F̀�	���Y55gVq�u�(����+�&D��z�9�-7l�ukf�3���RI�&�B2)y�u���Mm�l�1õͯ�2Jֹ1s����/��uŷ3v}��f�j��*/C7������ؠ�&�׭���ws�l�&<�ߤ��w���r��M�1c�0f��:�`ɺ	��'�|��"�&<F/?9�w��j����`�j�Qss+:ܬ���{+/�0�-L�nfB-�j��E����~X�e�`�DGfԲ�t&ù$nЈ	W4��=I�\������dΥ�����ل�u]�)�^����3䌭u[�9�F21�:��.�c^Mĺ�>h؜�^�p���B��p�BZ���!7���N�Eg��9�'��P]H��M,�K���F��f��9��lM���,Ñ���'nV������wS�p9�9�����[D+P�!퀄���,Ě-�r����\q1j�%����s5��pfe��R�[��rx�_�-����C+��>fԄ�n]�j��&ο���|���0��܈��)E���� T�~y�$�����B f�՜b�<�B�j�j���+�@
g�EhfB�Ქ��Л[p�h2����*n�;7إEW�M��]��s�[n�$��H�z��J%9���dR��H����6�md���5]Fɺ��-׍_0�odf)oh�٘	S�S���U��fq���?�'6hĸIAb�Vy��l�S��M/^7�O1Z�8�I9f�F��3p�T���&<n��f���dЄ�h7��AwY�)1aJO�m眚�[��f��,�[y���n����C���PMҿu�9��9cv7FMtdF-[N[��sIb1�C�f_�'��+���d&�f��uj��ل�u]�)��b���3䌭u[�9�F21�ڼ��^�Ǽ��u9�Yz~oxY�	S�R��rp
�.��P�9�&	���^�p�,�C|!��"i��&�%xGB��p�얯�e�i4a�C�GB2��8���#f�M����s8��o�W�v@BSe~�b�X9����(��W&!�������Ƃ��acfe��5<(�)���E7d%3�V(��}i�Q��u��m6�&ƿu��.G�R3֪q#&:�qBj;P�PA��	��u��� �0h��)�̓-�ˡ6���_�+�,�f���r������YlpZ�-�erܭ�U�Z�M�?8o��O��u�ve�-�+�)y�[�d��S�0#i��kX�s\�Sp��ߡ���Yb�T2_��(�������y]�����	��u5hV}]'{8`4�ѻ�8�L�OhN�5]}6fc&,���34�*��Mx|����}#�%����j� �pR�ub�a�ƺ�q7'��x݂%L8��eaM8��&�Ԙ�K�L�Ѯ_��Q#���q��,9a���W��FjLj7O��!�ˢ^j��7n�K��4�J�י�^j�;��/5��ꇕ��MX�Ѯ��ь�H���AVjɄ�O�lB�hĄ5�p9�ᘙj0˼m6��5wsoĠI��h��"�ær���g�ـI0r����O~4�n�.���ڭ�uS�X��X7��fY��3jjb��¸���D�X�};�N�Sn����_w6������9,��'`2�����p&2�W�j��61֩9f��k��a����f6�1��y g��)h8]Wr�.�kc�Ɨ��#���
4s�\��-'�N��_����/b]�o�Z��j�T�GO�� �=���߸�_�Q1a���l6t�ԘI��nw W��2��p�4p�m�	��S1`b���g7���S8��W8��h#�r|��y"��,�f#n���n��!�f���f���
[�K &�d���q��F�
��s��A��x�/���a��G�[�ǣ��-DjظI�g#�5�8����Q���L�g�.o5k'b]
�`�CגE��Lxҟ��f�����[�[jfq������2hΒ�p6��<>x=c������AS�;����sm䰁#&�s�u�^���r��p��@��ڑaS��F��j��$���g%WW���,���������I��j�{f��Lu����w:F�(u�Q� �a&A6R����5��q,^��Β_=5�Dh�Λ��@�I��y��Ѫ�O��s�Af��A��Q8p�8-N�c��)��v�����&Y@ЈR0\���2�:��m��&6��2+��@��df����rVt���Sq�����iX(v��`�b�n���;�����I�7uj������8�M-�c{ᔓ�26�:7����U�f�6���=���_�k�&b]��*�5�[L�ү��ؠY��+��9^�l�nиI���/~2M����y�f��X'�\X�Y��q���r�g�7)��Kҍ4�`*�h+�l｛c��V�X��]>n6�f�[NL�7�Hl^ĺ�6`F�%d��<�89`6�$e�o\]�/VFL���<51rn�����v���beor2�z�Y�p��Qs�5}�ꑁ#L����R��pnY������kN���^��OĲ��B7`FS7�I~Z����p�,����C�0I�mn<6Ոi�V��#�f^M4a�SC��_��^7I٣ԙ��ȹ�jظI�_~G�^�v�ݨ�-�L�d*������.��ܐ4n̄)���Q��ھQM�]��uQ.�ǐL�j�Ӻ�9K
��Y!j޳zj�1mK@��-���I���\8b�8[�����@���ڇF4K�4�:7Km=�L51�^��.���f��V��Z����O��vs����#S]>g�l�Nǩ�nAX�o0�f�F�33�Y��T�Xf��'�%�zj
���sT�@�I �y��Ѫ�Onn�0���$��Ɓu>L�"N�@mJ*H�<a�� � �e-#�����AS�؜vf�gG��bf���[���T��L��rZs7gT�B�{�7z7�,�{æ��Y� �MJ��[�SR��GS��b���)'5�eKma�f�������`Ԭ�&R �����3n"�e�]�!��z�
Sz4G�6hV�h���c�6���d����e:i�45�{i�W@��n��rS��xn���C)������?8bܬ4�e��]�ؗ�f/���1^���e�>��r�^��-'�n����9LMĺ��̨���T�GOێ�-�EY�WW��Հ�:1O�F��[�&Er��]8p[��MN��+x8j�]��� ��pĀ��^*`v��-˵�p��Z�ȿ,�*���'bY��g�0���0%?@�׵:\5�Ũ9�6{HY.I���,p�OL�Ш�B97�j�	S�2'��|��I��n�y5r.�6n���?��i�W͍�Ͱ�fb�;�������.i3h��m��Lxғ�#f`��S�Q�uWja=��]Mɚ���,) g��y��y���������w��#�(?����\l��RO}䐉�1j6�ė"6��n�z��j���j�n�]�heٯ�d9�4`����I��挻�+G��|�l�D�R���!�̇�f���Huf�>؁"���s��Y򫧦����Q-�E����Ue��\�{h�,8h8
b��	S���"Pہ�
�/O�dmZ�z�����>�6hj��nq��Ə1��	.��
Ss�]�[.�j��{,n���&۽�`��6"+
M��M����27'Lu���@"g��I�.g���Bs˛��i�ei�̺/Lb�ufVo�>?ַ��9ۗ�Z�I�'��KcK��5� �ILf/d��<nw�l^�s�A���Uݺܷ���]U4'��F�[x�i!8�5�V���u2�^���,0L�
��\Ԅ�a�[Ӆ&��V�a�1�e�KL8�:7h��	â�a����^�0�Y86u�(&���rpb�.+'�{�F�˰huQ�.�^&�Mx���>�E36*�&��p2�U�^�M���2,���e�5!�09Z���]A#Mۼ��E]Lp���nmT��a���H`؄J��jج��s9!��[�})�Y6���[�3��̦eZ���r��*Y�o�2�9��T��*�t�ׁ̧As_���eg�\�eL&-�er&�ɸnp�D�ˆ����E#��==3W����P��9U�<�B��)�7��-�G��j#���[�s��4Z��da�8Ts�Y��:ί�z��㊆	��Bc&��w�j͑���ץ�Y�{r؀YG9p�8�XȎ|3�n�E|����@�e��m��ӥ���\���ɺҚ�|d�0��ss�<9��C�5f��<�,���@����L����^�7�)|��z��6;��+���~A��Ë��oȿ��ty��@�����@���X'��^8`�D��~ml�t�Φ��#����\�'�2*�>��1�{�#����f3d��R�@6r�����J�Df��cE̺�9�b��l���E�K��ZfKf���w�.�;'Mס�sέ��5g�)2C��pu��25�+�v1T^�i'���P_�h�,v7�MN2������U��
{�#FN!�"N�@mJ*H�<a�d�ש0��:/tl.��]�W�6=��Ί���m���W��j��-��k}�`�YC2d�_v��i��� q ��C�M��������;}��xcj܄�n]�c��Դ�pV�����xʯשY��B�FN���'��7�|{�ƫ�uC�*m�J��dhz�ibF�@��X�}s����)�GL�ղ<�O�B�+�LSQMx����l�[
n�B�/s���>b|�Wp�u}��M�������8�~�t�H�d�4A����P�.F�5����hN_�r栽A6`�Q�0�����ſ��n�E|Π���D�aa9/�l��j��UZ�����\�k	7���3��H�,^�5^��6f�7� {��A�:7�	�4�)|s�Z2d���:�9��m6X��y���O���u���e�� ʦ��r+Ѝ�u_ȓ��1�rË�MĪ��R��A4p6� E�KY}�,��B�#zcK�t�AH���0~��F&�_���� �Ɵ�1�^��e��9'öz���gs�-b]
ǖ2Kf����v�]�%,Mס�sέ��5gé�	�Yz.��ej�Wj�bTss���J��j�rD��l�gr��go�qs�j4+�я9�D�8!�(A� ��I��^�>�,o0K�J��\�۠�M���b�+l��73��,ǅa��-��밢��N��y.&���`^q� ��Rw�c�)7�_PS��K�̹���Q�&\u���l�OMkg����{������M����©ܞ�dt�o�;|��cRMC�*�9/v�8��)s�X������z����#���ͅ��.e9�0�kA'�TT��}3`�,�햂��_�eb��q�G�O�8�`��qӬ=(nz!]�w �/9`Ԝv��d�4A����P�.���.g�s������Y�٬�
������B��՘�uۢ��땬c�f9/�l��j��UZ����{��~Y�Y�����`��o�±Nkc����+H�ݾ�1�]*E3�h
���V�D��1u��Ki����`��Qc�u:�؜gl�T�Wn�Q��y�u�*fYnxq��X��Z�r6�Φ��u)�7�fQ��p�j�C0���C�u'�a���L��Q�����@03.���u�s8�ő�ƪas�-b]J�c��%3�S��߬����WXס�s�m�̚���ԝ8K�E2�LM��J�]�7�`���e���Xl���C2���э��Z����G��B"E���� T�~y�$���.`�,�+���wq�իM���b�+l5k9�W��ke�n`�*Z��7�̍��Z��U&g%�"7+�L6l�'۲Z �\Y8m�Iu�\�p�4ɺ��i�":4��7j�h!�ƌ�0�_�7�ʘ�x�o�Qs���CW���Esu�~�����zѪ9�ǔwhV�����/[�Â.N����:�9�+��ҩ�f�{�&���;����SU�z}O�mR7I�#�����X^Iբ���˕s�٤0<�����͢�s��t��u��w0fR$�n�Vo8v�V�.�}9-���e��Mxү���s�9�u݁�ޚ^�$ǎ���Qs�u݊��6'�ʻI\�y~g�e�FN5��ؤ�gD�$x$��] �s،���lݲZ=7n�l�MA�r>@D�$��T��� �6$�ws���벼��nԬ$�[����������)��.����<�2_q9h1+um�hW��Qs<�I֙��7>�ٞMUo�_v���Q?J�}�z�~�ĀY��!�R���G�%����y��B�>Xl�Ǹ�f]H`Ψ��u�?7�e{!?l��G�ܺ�9��غ��u�8!�(A� ��I�U*� �e���������צ�G��k�q7KS�*���h��as$��9�,4ûb{��U&g%.�bc���u�2p߭@�ݨY�Ձ��ؤ[��
6g<5�p�|7s!�qSd��~i�9��,��W��hQ/M8n�uh��j63�U�_��bn�^L�#u5�<��j�����`y���;�Ɉ��b�T׷X#5[�34)\��*��g�j[��Z�f!u�z��͓9��l`yŨ��=���$�jTCs!.�YM#[�:g�;��ϱ5Z���z�Q�.��ƞ|n�gɻ	Sz4K��u�]�Z�f]����$9&g�����]�m.ؕw��O�Xu��]��ݣb#b�M������1s�Q3���##FNd����|H�t�Q�����!��R1���j��nԬ$�[	�T���͞S'b]f��p��9��A��p�E4p���J?4j��6�:7���F�6U�U~�J-�8�G��oWoQ����G���Ԇ�$���{�7��M��|��z�%�t��ݺ�>�*�#�e��7`f�k�.�ߜ����mHM�S�	��@	B�'L����P�.+��^H�G\N��6��}�7�f!�
f&����x�=Ǘ�fxWl�V��d��eYllR�-����pp߭@�ݨY��gI�I	��5��B��G�&b�R����*/c7E�����ڀ1s�V��hy/M8n�ub��,lf*���ܞ�d�+�f5�<��j�&�:,8qu7b��9�u[�YA[�34)\��Z�Y�e� �CU�^-q9�YH�$]�T�D�]fVby%U�Rw�>���e���Q��ɼ�N5�l1W蜹�`��/%7ñ�\!�2�/�ɷ"h���p�?���21뺻~�ͺ��C3ާ{�6΍�Qs�u݊��6�ʻ�!��',�
Y�G���º�I	�� ��s،���l��x�Rs�����Կ�uK�q׆Mې��ơ��Ǯ�j�5+��V�9��MSb��D�����S09h~@εa3�]�F��<��&�����1æ���/[��G�(u������r��,�n�q3C�8ҭۦ�7��M��|���͒�q��hn�UY�.���`�lW�ZE��7��,�b뮦�)��v�����&Y@n��>V���������צ�?�������f�L�t���=W���h�m���S��/�ѳ�jB���s ��m���T�׭��u3�][1�08���i�&k���򼻶b��b6�Np��!VL�nj��85�o�ߍ��6Bx�_��Z��[Y��5�O��&���ݰ�z�ɠ	��X�`Ā��q5r
�����F����|��4Aɰ	��]9h�<��',��;8f#GN��/э-��Ki����t��I�$R�u?�o
5j���V���pޮ�z�I�Y�r؈9B���([�u8s��pաAg	�9�ݐA#��� E!;��t�l���*�^����F^�M�[�[�132�I�gs�/���Mĺ�����?3�9aJ�݌����"�YꇴE�:�.4Ǫ����"e���Z��Qv�.9�2wM��ЀYP7�� &�g�C��Zw��y�@kL����r�4�s�ʹ[ؖ19��f�%��^��U�Y���9��9І���`����L�ҫYBr��5�/� s��,��	OٺM�6���ˢ�w��0�ue�&:GqBj;P�PA��	�, f�C`���rkx�<154�i�V�p+�@���ZNh4\X8��dh3`7b����'���k���Z4ϫ&D��z�9��l�upܸY6��PZ�q4.�{�LJƗ��ٽ��� �1b�;˄�2��[v�rc'5�oh���0��܀!��d�&V�ͭ� �P�9��br���ԭ�#���	���s�`Ā��q5rj���Jof��ox��{��aׯ��]g8O��Lx_D�v�Vjɒ���C�e�&��n�K�⹅n��	K�fW{�0j�$���������`��.GN��-�� ��W0Luh��YnNn7�]R>9j���H%;5`�Ȣ}��L/��y���S�bSl�tcfd&�d��zPV#���u�����g�#'L���U>��)BY�[�9��(B�ɶ�p��rb|�/�,6+��[�F�1e겑��-��&Luh�,�Kz�n܀�B3w���
�Ժ�uA#g�5&����@�j������.c8r��ݜ�N˫�#�0��0�y2�0q��=9�q !���¶vјaS8A�f�9(�Q��u��m1~ŗE��Ҁs�/@��FMt�(��v�����&Y@�r� ���33�n�Au4�i�V�p+�@���ZN�-w1��̀Yp܈9N���ֺ��p�u4ϫ&D��z�9��lb�V�ܟ��R�h\������/[��{�EX�Č1Ýe�f��$����:�ب�X�};P�3�l+2�I�����<�a���Gǀ7)(O�a��Є���A��U�ƗNMx])3�M���~u�9�Ȱ	��Kb��A�)ؘ	��l��۶RK���0�_t�z�¹����xn�9p�RuSNq5Ib�""i,�3�9�ˑ"e�}9��3�
W4p������y��8=|.+�7��Z�Y�Ó�d�u;�O�S��(�ҍ���L2������I�.e�<mN;1r���|�)BYj[�9��(��d[��s���S|Yd�,����5n��Qv�����0ա#�<_�ܸ�dg�C��Zw�.�b��Ƥw�f�D`А��Y�-�ltÑ�Lof�W�:-�B���؄�ÿ8b��
	'��M>��L�ҫ���Ec�M���Ef��1�&<e�6E�\����"��mЬ��ue�&:GqBj;P�PA��	��u;��X]0Ͼ�whu̜pr�e2P&fU�2 fvE��H����1qu7qv-����وaS�y�sn�|Z�	u[�9����I�������Z��S�d�1>�,��Ss8�Ͱ�e��͢[�]9I��,���4?��Lݍ9�?���_��0Wm)��vC]�������D��z���j ؄�����Z��p�d�M�0���\o�7u�^��LFN"}��ͨgX�:2�،4:4��yy�.��,&�߀�Ɩ�Z�i��c�.��N�nm�9�,���ֱ�����^(шI��n�����#����<[d��A�r1�:bb\�R���h�\ p�$R3L\n'��ܸ��+y�Lƴ��%:+V��'�����-��w�9�Ô~Y���h�T��IN�M�Iԙ�$���1F���fPr�X9h�֙9���Y�=U��<���M�@��j>��������oVj�j����e����|���<R��Q��t�-&71 ��z�`�Ĩs�2�!S�hf�Wvۭՠ�ᯙk*�Y�D�+����嵕��ɋ�%�L��%tH��n���:1����M�2u[�Y�rb�$�q�leܜKn�up��pNr&
v�lj��xxd3p�-[��2Z6EX����溉1<�n�h�,&8h�'�$=��_8��"s8���',6�E�6F�ˈX�hn򙱒r�N�����
���r)�y��,�e5�������̢8i�R��җC�̅x]�nG(����t?��$K�Shη���B�z��5�*��
��7�2_��@�N�ދZ��9�O���j�S�	��@	B�'L����}��r�+nV�)��8�=7\�a����r����K���L�%�L�����I�|��%q��A*u�iPq�V���yw(@s �#S��/�dΗ$��	�˲n�����,�[&�-M������5��B���Z�r5��pӅ�r�h�t��+hVo$�H���m��̜�r����r�XWp�P9õ�G3unbA��l �D���b�5�Rw��)�%p#ڿ�)��	&�48lܬ��fĈ��l�xX6I2H�/��z��[8��ɜ�b�$}�@�huQ��M��x���<7S� �Y�5[�l�.-㥠f��r�T�.e6pÁ*Ygf��y�W©h�p7�fl�I��r�\��ok+f-ќ��,�$E���w��`��ߖ��ݑc}"ו�fn�Fܜ?~[&��73��$q�na�j�U�`?�_�:5�
0d�11��Y�<��\�J6כ�p�L�:�F4p�\ٵ��?ds���$����n��+R�lf�݌�+�Lo怵�7p��TH9X�9�V�@c�*���v���� ���N�z��p�����.+��o��G�;�nr	,�+#��%xf10{���K�vׁ�s88fv6I���X���ZlHG1�I֭0f6y�oz�:0�׍́v�JLxү�#h�.�Z����$�_���6�jݩ'f���Z�I֝^l���}G�����<��h��t?�Gx������3�fVYͪ�G׭�b]��_�l�$��/�g���Z���r���v�+�� �]�X����xX����H��NW���1S��Ǘ�������Xaos���(Ud��v[�d�5ƍ��AS�vavs��9�$A���>��G�.�]917vmĄ'��?��65n���S��tx���$��u�~5ظq��O���)�f]͸�İT�it�s�`��]w�����+	-K��� ^�WG��r��C���tO�S吹�p����tu.`b��n� ��Y�I�#խ�=����&P��A��j�����/�Ϋ��ň��#�"s�G�K�gs�/��d7�I���Y�۝�h�����| X�b�"N�@mJ*H�<a�dU6����-��b�M8�g�Wac��t� 35�
�Kj����V���Z��wh�&��ͬ��9+�K�;�2�Ug?a�����+���h����̀�Һ�o��]J��3��ε-�\��<�>J��23�1�&<�ـ9P��bZ�b�T�s0]2��C���l���8�f�ޢ��A�	�ȐY�D��� �,ؼ7bYI~W���%�rK�Lx�ߛ��0r!�S-;��K�:5>0�c�b�Rҿ(ud��9�VnE�$	���,�/y9�]���\hnN]4I���]0nn)�J��8no5�$L��R[)7&'<$Zo9n��`sQ��:5��f_	g��ٜd���S�Z��-���$k#�}��d���a��+Jٲڜ��21��ϋ��^�՜:233�h&�'�	q*m�-9�0�J�I�G�C�[��Z����&���d�F2�T9�R���{yyͰ	O��y�WV��^�]ga���v���[4�
��{��S�Z~�����I�F�s�3�\2C����Ј��v@S�Tm}��7nhyWjG1��1U�ĻYY��f�ڍ���!E�:3�vd.K�L�٠A�fp>��_�er�\����S�V��P��;�.���p�M�҃9m�#��㦸/fV����a�:4�*��&ƿ(u��s�2`�Đ�7'�3f6��[vl���N1�	��q8�/�h"�e����haJ��n���f�h�$Y��Vw��ϻ�krSnɣ�A��/J���Y�6vP��Rrcf|}* -�#��a�1Ư)��]�j*�"�%X/���\�%	'<�7�f��n�Ꟛq�6z�L>R��{o�8H�?J��u�?cX�f�6��ΆZ�빑u8cY����nИ�X��~�d̈i�	S��_�sd�vs�S�qBj;P�PA��	�, Ë>�pY1��fjܘA#����`�#���E��9�.�����xB���&��QꎣK�Xo}��j����t�ڛQ3����d�EZ�5ZP7fMĺ���r���1��7���/F���+:��$�v��YH؜6b�4n�\(���|0N�]���OM��lܬ��x2ɺM?�覢C��m5��,3	�N�[�,6P`��\�����q;B�}�s\��5�I��������qs;�p9]�*ws��H�ݒ�-5pĀQ�������嘁�(�[x�o��^4�,8]����vu�p2؈9�o�A0����l%Ό5�(�$H��>�+��Ӭ>ʗ��u>�����1��b6r�Ĥn�50�:l*i���a���OQʮۥ[�'��$}�,|ɲXʷ���gZ��'�.$5��R_u2d"�e�lb!����UN���G8͍��в0jΛ�+Yw��+|�ы���uU���')w���O�t�������e7�=��l&���7�I�p4)���}O���99c�6[VD(��]ȶ[��6�I�3j~Y�����"N�@mJ*H�<a��i4C�`��Y��c��an�U8��A`c;��l ��X��!6�|�m���/��~����Jn�˴�!R�B�������I�?���q�FN�v����sq���֍���u3\�e�F�r��1��&6�J;5b���.HpȜn�$R/f7�SR�j�����
9�$����X|`�b&�ַf1-8��c��6@�u���\��d�F�؍.󃽛��T��+�s����f�/Z2b$��M��f�خZ�q�~151Fo��l,�Κ�as��9��>E�G��(�Vz�Vs1�y.w5hZ�뿖h�.t1I�8����\�[v��9	�ld�[&�yy�z׭�^d֍LҘ�]��Aw��VT�0���h�b��]����[Tr̄#��<��<R���"5b&�B\�{��Ś��q�4�@��G�"8L7T/9r���w$�_R1h�����#���h�,χ"s��\XR/��v�^t��2p-GF6[�	W�i��n��$�����	�������H��5��5�J��!=��8[-4��t,H[�ef����r��?�}K�LxH��<WfU�O�1]w�]0/1I[գ�4[�K�ӟ�����!�dm��kq�13 ��/Jݍۤ������f9`nہt��D2'ܡ��8��ܢ���ed��	���$��֯a��ėӆ/�ek�4Y�Gh�nYr��s�Lĺ�4w� �Rd��	O�S��7��:�:4b6s��9��[e8l.X2�Mu_�A�<Y`�1��(up�,�kf+�dy�:7����s��P�͡�uX��Z�.f	���ͧ yt��$�l�vpԬ��R��5�����5ᗚ�S��p�b�T��As&����6���HuPܬ�1�\Р��&L���@9T��ڒ	C�shbs����"��i��1s�Đ���8�Z2d�N͑J.�fb �zbs�͸�X���H���33@�&<�#q���+|ё#F��$kќ�r�58b���$y9�hb���s����s.�cP���FM��e_�f�h�X���S�&ZY��d��k)�	O���m�3�).�Q3Z�dĄ�n<9W�Lm��n��Hf���*^pO�fa]�Zwz�7���Y��j�\χ�u	�.��E�Mx�G�37��̦�ܱZ��"Pہ�
�/O�dA�f��Q fm.�i�\�g�sNol���,3@���[�y���s����r��as�-8p���9<��fV��:edqk9��m�ed5���ה�Y�7��a��kt�/x�l�֚�ѵ95�O���f�y�l��E++�����FΘ��s_�g�=m����C��0��H�s��'J�F�aƍ9��n~��#k]Ǌ�i=�|��j���9VЌ
r�S��6d�V�~'}Z38�!����qzM����"+�M2�6r������a���p�s&�j�Օ=&ֶ�67���fƨ00m�a��uu�eaZ׵>=����j!$�t�\8K�Mҟe�`I�Y��'Ί���˕��>�����~�.�R?�q3ed���z�&	\���	}�]96���d��h�sɈ	K�sG�)�եowW��w0�*���
��'�,sSv�-��|�$�\����}y�wW�̹4Ϛ��q7t^���vS밲�:-sx<iŐ1SE?8-�{���%���kw ���]�y&g������(TS5�/���.2��&<i[�-Չ=n^�\��6�f��[|OV���?�S����@3HR�L͆����V��.g3��2H��Y���9hE+�>-���Q�4+��Q��Ńf���ȑ���Y��In��Y@�#F�$��ו�<�ʻ9�.Q4]v,���r��;���heي��fXBf +,�����!*9/[���`�;B��5��p�>E({�9��<�C7'��3�pg�ؘqss�l�R'��Y����j�ȉV��'G�B���8<���\Xw7nд��䦗�4j�
�8!�(A� ��I���h`N�c~���Ay!?�J�p!��
�}-j�E�nn�z4��q�n���\k3IbE(;plr��ꛒ�sٻy�!F�@ں�
��o�F��M������ S���Ӻ]����K�%D�DdZ��:�wO�c6Y��Wa}����Ŷ������d�9c�a���mq`Z�K����,6_�Uf㦉�l���i����6o��ڸ9�ʳ`f7��d�e���<�I�'���s#o��BFM��co����
��C��k<�N���`d������(B��j.1���F3u˙��Z�)[��G�\�lK���xӫG�oyn�s�ܸI�4r��/�w<:մĨ�!rn^G��y�92�[�8q�e��M���纩�HI�b������_'i�������ϱ`�-�,ڛ�w�-o5�y�`�D+����a���f3�I}�n�����0�@nf�Z��$˞w!Y��X�"�܍ssޢ	C�h�4ܜ�k�MR�e����0a&Ƨ.4��C%����nΚ� g�9��K�&ZYV�f<�cAO�XV\���f����R��"Pہ�
�/O�dY1 � ��y�4��Hr�,�ljӹ}�"s�.�ű0���C�� f�q�N"1�Сnl���#[�ٕj���jN�]�@�-E���,k0g�"]�Z��p�L��!&5�~�bN��~�:1�cl��)�_w�#sn�}�n٠A3�z�3��άE��`.p7Q�����f�]	8j؄'��xխ����;N���L
/[���*���i����5a*[��y}��oc�D.[rnǪ���*��"��������V�abbꆈ�8��`&j�L�mV��5b�,��ќ�pvh���G&���� ��t��tݥ���	�bdb�[7���GS��^ì}2f�S�:9f6�0{�wz0Wj��q�����:�S�{����Ac���f$8V�
톯 8�dL��T#f�v�5���Seoy��ޱw�SĺL�� �@t٫�aH��~&
�j���v�Y�ШI�w��#����]��z�8>@��Q�V�JW�0�?�mލ���J$�|��l�m�֡�i�\�e�&����+�8$#�e��9�<�R�N8���\�˝+�:� 8E~E���� T�~y�$��0K� ������f�e�iy^�`��|i,h@�t��۴1U������$m�R�|��5���Wϻ//3��	d�9�oԑ@F�����h�|Vy`\MxҫYO7G:4S�~��&,7d�S� ���bi=\���r��J�����u�0sГ�������rk��$�;����dn1��������n���{����~�7��e0�d�v,�3�DVSq} s���r�$ꢰ|骹��ߍ6c^��̚.�.��(��@�s� �n���VjY�A�D��7	��5���t���^���u���l p��=2`�R������S�w9�m�0պ0�-�s5p���V��(uົYJ�[��$�3��@|.�٪��̺�.,*7qƯ���5r"�e�/��Z�`NLx�G���yŶ*�+��v�����&Y@Ƞ� ���箜�9rքMmZ`V���s�3S���M�1f]^b*H��Z�Y��0I��Z�+�h\���]�b>�b���Θ3m���}��Y5�p�$��{ݗ��[ͷ.[x�n�\��<k�F�7ǩ6n6-�h[��Tf#աY�`�,1wDL¢(u'�[�,�[G&��K|�̨1S��� ��ɺ3d]7��������s`��,C�h��ehu���]fl�BYb`����u���Ky	��:���#��D�Kl���.�\�u%s�+H��a�4B8p�ԌPFf=L1��5Iˮ(�M�>�^Lx�n�v��4$�&b]���od��zW��l��8K�3f�uj�Y��k{1��κ�ޏA&\eh�{+�%���rs�����lr4�,97���"3pa�����B�С�'�M���Mx��)�,��N��
�!P�Q��V�(3�g.[n܍�C��"P2r6�М�'|v-Z����N���c#�8كsp[��[��͍5X<r�ul���e�q4b�ak���|��)m���>-��t9�)@ �5Z �۔�c����ByH7�+p�+��{LDO!�W��]�c���v#'Y�&���M��77x��4��Pwe��e~�I�2b�u_1dn.� o���3����0�����0�%���Y.Wu�ݜQ��cs��\����~ݲ�k�(ݠ��f�f���'������]���u�db�4���lذ9��)6�`['�$PC�̂ ���uf�,;2��`����l~�W���4��|j�Y5�dhȈ��Q�z	��<�ޅK�֝�b�q7�&Y�,��Q[��|Y���V5n�|w�����.�uj >I6}r������qkVr��D��|_�]��}��Q��g�&���jY�i�̴�`�1I�T�Wn��j��G�#sB-�{m�4L���
>R��y�u〛�����Q��ﱙ��ȉX���46$�F�6aJ�>4�����T�N73��"2`�$���Y���ֱi��9�$�N�9g��æ���"Pہ�
�/O�dY�u�0`��R4s03D�&9b��$�3�}fjp5n{���ȩ|3���	��r�|�R�|��"\���c��^�l�4%&<�uj2wi��	H�Y��V���%=���[5f*�&�
���&��ԝ �q�n�8	��ԑ�s.�͉Y�b�[>rn�r�U���ꢕ3���+s���/�Ƌq#�~]�M��S�~�_=7r"��Ѩ�#��5l��?�I���Н?C�T��ofA]��I�E`����Y��xC����X��f��f��� -������ƛr��$�^N'�S,"6���8��RL��Y%0K`�"���L������}ք'���9������������Z�l��48j��i��+B�������Y6p�����[��}cea$�Y�7q���Q�\VNĺ,�U'�񥶒h<
g�����qBj;P�PA��	�, ��0\��9d.����,G���6DW�i�,�e{�0SC_5l��e�L�p����[�-�$m^�E���p�ՄJ�2���7�$D�b�Ą�n]���������/�Ną���~����huQ�e�M�����"��+L�ڰ1��8�r V�.LE�R�$7�����ӯp7��C�2ۓ�|��s���"����#։)ufԨY0����'��M�9d�q������YS8벀� \�W}e�����&Le�y�͝w�z������M��IO�\۽��+f�n΁��,3ɺ��E%g
��TZ��/�w&}[9���ZG5jj�8{l�,�9�|y��p�]�����G��w��m߭�3 9u�O�8Ĥ �����d��pĴ�k{�_�}�%�?�]�^u}h���21���HuS�6/�̙p� Sw��,�k�FM�{E�s3hNC7I�N��jl���K���mY3%}��EiF�m�zGYu]� 6f�����z����Tsb�9�Ib��Zٵ��K�ʿ0��J�A#'��#y���u^�,�U_V��J�y}�,��Ď\��/�e��k��	��X�Ą�N�kn��a&�~7��s֮{�����Q#���.Nf]6�:|�-�������L�C'7r�Ժ�Es��ٱ�L?@���f�f�3�����mL�Q���]���F�11T�R�
��C�i�+8���y��T����.,+�&��G�f)�Y�V$b]8��N'D��%�_�0�2l�c������q9��rfS��hVr�C��C��zaXN`s��n=3���$ܘ��؊�lB��9܈1���8���W��(ƬOt�B�f��nض{}�<���1�G�[�o���z�`�$�z�?ۭ�2۴�e�怃��FN��Bpv=�D�+�-\�⺘ÆM��Q�Nr�t��T_\kS���u�&^�~�[�#/Ywy��͂����k��;���Tm~��,3�W��/����$���q�s �L���~��Tfb�G�[�'���<
O�u��h��N���̽��`�}�Ng5�Z�F`1�Usv.��NĲ�ף��z݊�	Or3O(�n��+�u�ǁZ��33Q�f�_d̘���ll���������.ۡ) �*�;��p�܏��Mmr��K�sj��x������e��[	'��ub�̛���yݰ��Ӹ��*-Tl�l4�����6b�Dĺ��Ano!�ȇ���5s ~�¡���;P��$IN�ey]����]����1�)��Vn�n��J�_v�s�T�Iy�c��:�5��@�s�9�c�Y�u���4�_�C����3������#��K���N'D��%�_�0���}��I�B��:�����4�>��]%7+��gsb�AG��s��/��LN�}��+�F?��5N���,yꖗ�)5s��΍7G�}Oʒ���<�2^ȪlϲN���j�:5���֢a�.�7P��1��aH��u����J�"ts#�hy�r\�j,�r�zK�v������]�Έل��,:6j��d�{Yށe��0�n��i� rb\_�n�#f���fƒq���oȾ�N���D�+���a�_�nԄ'�*��06dfj��,97���ՉY��GK�9J�}٨�ͦ�$�tp��'�����2!�'8I���F�\a9f�ej�ρ���3Kyu/t7�R��/��&��p�z�ev������ou���^��d�,�h�&�u��K����&Lu+�>�RG�[���J��XФ�~��F�P�N/1�@�Rb��Zn F=5���x���eY51fpVJ�p%Z���R�]�3����4�$����o@ͱ�L4/�=�P��b0��u�V�T��H6�un䜺+��i�&��S�d9KGN��9qI���ᅄ��p��.�w��j�5n~�#s��ac���z��i4I�E�;��x<S��������M������
���YVn��9�b�_4��9�Ki}����Q8���-�`n��R��"Pہ�
�/O�d�vb�X��|4��A� ��hj��12l���/f�63��p���.���g��Y�`��J,�T�׍tj���k	-%1��Č�d�C3�a�����`f����k�r{�s�ݺ��ޚ��M��f6��"�u����4h�D�+��p9`��u�I�.bȜPl�,s9տ���Qa�ۿh��4I��-.4lց��ۆ&e���g���F�֭����2��&�}7h���"����u�z���	��Kc�Β�x]�f3��zb�:��q�S�Z/0f,'A�U��>n*��g��@V4�m4d�8�ϛ��۸9u��-�B�ĺ��$��/��*����&��|P6'�t���v1��F�9�&�#'9n��4L�!s��k�Ѥۛs3�j�Cĺ��{����s8L����!aaj�����¿FfbꆷK�́�LM��.���h%��A㹫�/��ݜ�j%ݏ �ۯҚl-g =ƺ���z.W׹9A�Ѳڍq_��~<�͌����]��̋�T��P�Y��΁m�ʨu)��k�ܸ�a\��5�u5�&.#ԡ�aW���q�'��R�Poj���Py��Y��%�Lh-5�m�7�&�إ�l�\�heY(�z��w�0�^�`��y��{-;12�0q�sj+'n��r�9<$����hc�{ⲩ@�f�������Y���FN���z��9��ܠ	K�e�q77\�B��]���Z�3k�cX�n�[ge͜IY#�-T�ȕP��d��o��c��� �9l���1C�5^�f�D+K�>��^���&sF-��9���_�k�.K��)��v�����&Y@�vkw��~f�L5HӴ�.υ����t倘��n�,��.������l�G6"G�����~�.hk*ufn/�!&��{�N3P2�q(ԑY��E�fԸIE�f]��(r�	A��X9��導Уk��G{�P�[�hogy'��W'&,u?7%�Xa��a�/�u��ſ0�k�B�o+l���uJ��v6p6�z+:P�&D��,��H��q��{�4r�Z�dj�Z��f;0)��� �J1p�Kտs`a���2f��C#f�hଳ�aS����F�����0%_��ٴ��9Ų����ń��b߬�/p��E�������A�9�ԄH�)������e�:3��z�Y��y��6f��t���g3:�Yff�ulĸY3�LL�v����ѳ�麪aC&L�ݬ��s���)��Z7M݄�l�$��	���ׅr" (̐�b!9�{^^��}}�s���aem�p�v7��D�s��T�<WN̺�y��[7��I�]�U��5^8h�S�s�Nυ�Mh��>�W�pvg���N�\5j�I2�Au�ã��#�,�^�n�⊠#&<�����o����-��j���IwO��t�eSY�B���S���I�?��e�hbJ�a��r����A5��y������d���m3�®{�
�P�L�$��/��=a%����:V����z�)�ŗ�,]�輦w�-9�?|,�l�Q��b,&9n�0��oͅ�"��R��s�VLR�(u���B�h��s���G�S3�^��61����`�۫iz����~����ڭ#�z�=��u)��,�j�!#<�����Z�`���{�;�$�"��T�Y�5sԇ�nY�6���H�Mf���9����S�I0I�;vVa�Vg�j��y��J��k}�/+3l�w���ܳ�;0�$����jU���X��R��ܠ	S��f�qW
K�e���jŀ�&7�rkt�S�N��gy-χ�I?������DVI'D��%�_�0��Ni��;�Ќ�b.P2��
�M+}�M��Hg��63�q�֯2�d^������2_�/�UT5����fCbb��8,��ȩ��4!��%a����E��5=�5�3p�j�u��`��-���WsWMR�u���;_�֭*��u�ߐ�����/�`Ȅ�o��K��gxx���m��Lؒ�I��>+ǆMUM��k���M��bΩLV8c����N
m�Wquo��S��4]�p��118]x�,���F����8��wM��0�m~i��MI�"�-�]i1��#$Lu��zw�Z������ᆌ�C��Vo��er`9����ٜ�Kn�4��m��F71��9 ��r.*�p�]�c�<SS�3�����M������vM��E��rېqSw�md�1�nѸ9�^lb�?|^1+U�M]��YAw(���ғ�ߓԺ���#�9%��'0�ĕ&��@�ʭ吉A�Aw�y=6�2�mvc��Yi1�I��9���E]�_亮9+���z��������L�G�[/8pn�i.&	�'�af�/����BqI�\16I��[ͥX�'�:1p��U�s�� ��Y�C��t�ѽf��|�᜛3���J�E��)�u�7%g���©��+%����&����٠�#�B�ad#˂�F��E�;��ϕ'�}�7���u	�a󶩻%r��2�X�+p�x=6�����J���Cz7Õ%|����-���L�@�Ƈ64�n��z���âڂ~5��;7Ϙ���M��<��o�rl��pb_��.�U�S�[N��QP���p�耺���<��vs�d��^=5S�U���2[�c=F�M���/�s�����\���Ť�Pw�����"��(u`��p��0�>�u�V��m�d��Qo�d�lpmԬ���u�?6jn�R�#'�Y��jN�Qz}*��7�� �L��h���C����(u����Z���)�S�	��@	B�'L�ֵ��cm��if=w����=pԀ�d�]��L`6\�<����� Q��uy���#EO���VsP=A�	M�j�^�`6vT��P�Z0���z��$�Dwr��9�_v��� u]�z�3d���#��z����1j�$���ل�1���ʙ25K��8�>4&}�P���o��x�X�F�6bΛ�e|�����҅-��.��vA�i��ǌ3/Z�ɈI��9�7�|/��ʟ(�Gz�_Jd.��*��S�-1�"��"v]��*�˦�\��n�#p��neG���Z2���j���$��,��&a��3г�N7S��x6Oz��U�l�R�90D*�>���8����v��ޞ[�۷�hn��]n�$��_3��v�V�l�?��^v�nt�VN����j.�e�Χ"3��ǧ��9m�4���hN�M�Qc���9�Ux�j]>��$嗏�� gѐ9ݣ�e.���s��LĲ�z�=�ܜ!q�@�0M��e�6��Ca§(e[�-P��uJ�G��%�>0b�4l�q󎭖)2l�>����=�wcŊÁ��/��S��o��L���%n�Y�jЄ%�1��p��2n�U9�I��p�$�ޣ��Z2�����ޙI"%�
��|�YM����x�KX�?�cǕ8dЌ���qt����:,2G�2Ѫ2�p9{���h؄%�2�@�w��Q٬�U5�fM�ĸ����ٴ�80������7��$&uu،f�NJ8j�<���d�K-8#��πķ�!'i�����%1V,���r�����`�2+%FN��쏘������Š	K��p�f@�1v����M��j��٬��|�O�?��N��}v#�M��ky�������ȹ�jb�03	�l�xR�&ZY6J�
Z(.���A���|X���s�Cj
�qBj;P�PA��	��M��� ���X���hZ�/���J�_O���a���嶀��0� !���s��&�dvd԰�S����R���Dt�Of��Jr.�?2ɲ�ss��y0�}���ӊ^�Mm�9�20��́�MH�E72�O!PvFnif0�&��W�	CUt"�|���z��6pU��1+h��Lt��g5C�8:2r�����(��n,�M�Yj�$7�)Zpଌ8��I�5]�S�&Kg�B��7��U s0�����zd��1�29�|ױ���$�Y?3wo�,�{=e� ����&��5�c���܂�ZP�cەb���¼y7�!�GL�ٱ*�h��]�UN&�{wI���l��y01~��b3�z��eş�|on 7{�I�����j.���]җ�._��26��g�F��i�����7i�
���xGT��dVJΣ�AS&�䁳Ԏ6���n瑚.'ɨ�m�uO�<a����c\�s,^���U+l�^�ݛ!&F�5�Ȇ؜�r��en.�%E榮�K��*�nN�v��[0G0ɪE}׍�H܆���R_̄��#�ʱ��ز�����nl�$ɵ�$�9w���A����B��i3+`�.�c������̡��t��~��Ӻ�-�pc�u}���`����Kau�L�qmf9�84I.�1����r_����r�>���?���BB&r�"N�@mJ*H�<a�d}�����F��v�:�J��^�us$n ��	�§���l��2�2L^��{g���}��.�6W}�����'�4u+s_b7jj�cxi���"&��ul�wÌ�v���ȹ R����ʈ�ld�Q�j���2�#C&<��l}c�j��͑s��$�Wsܜx48��UPs�_��La,ӵY���u�	po�L�����>�h�n���լ1)5�x6g��/dM�f �I��)8���:��D�+���gK��Q�J�]9�9��v��a��-]�Iף�=�=$��	�"�������p����>���GL%�~f���	��<�z���Ϋ�u'�ٱ�/߸�������1�2���^bИ�X��~�`�<�7��k���T�9E�u��C��{U�j湯I��(u��\��q'	�N����6`�ĠY������<��}6\�V�]ͺ.,qTv��@�l''b]a3�r�b�����Ƃ�o�8���u��r��T0��ۘ�PW�&в&7M���Y��{����Ϋ���(u`[K�>^��Z`���	Nfɪi�����͓AK��= ݘ�Nĺ������ԥaJOf!g�̖=�S���f���[�Ir*R�f��5�ϐ�/J�u��j�h��/���\W~��)�z�ġ1�x9�FͶ�Mĺ,�Mܦ�!�Lx�G�1kg���aS襈"Pہ�
�/O�d9������x�3��/�n�YB�}cbz�7S_��^x�T�l�ln��I�%Jݺ�a�&7d��	��,�M,3�ˆ�� ����J�Q&�כg��������f�[ �,�uu���9��u[�j��_�+��I6\�6��l�XZ&����]rn�z�9�y�:8�|�0j�������V��z��܊��d�vS�f =�<J��S��
��p��T��Kqѥ�G��\�h40���)f=W�����1���j�����e��b��67��i�&<�Ɍ�fܬ�2��:3f�}k�faH��]�As�����?��X��$aݜ:j�v1h�e��uX�aia#`��2Y��H�;�g�Ь�?Ё)@�2`V��K.�M���u'��ż�0)}^���9	�����n�,����0b.�ڡq�.��L6�����ф'��GsƬ���h:�d��ɈI�}��_lv�Xc�]��x�+�&<u�L�!vhNL��m{)Ȭ��N�\�z�65gQ�i,Y���=6I�Zn.�}9�j"�e�6����e��QX��g�(9���8!�(A� ��I4b���B��x�Ը9�Vh�#6&f������A�*8n.����½y6�e��bZ�b�RFsu�H4C�;���Y/�$���8I��n����̹�dF��0w����;Ȉ�G�$�Wv#d��c%�D�+�-��8L~rC&<�7M�]Hמ��b�	������$�_td��e0�^ݿ����Y��u7s���(Ïu's�ԨY_���V��m�֑���ݰa#�L��쫹j�܌��M�&Ywɗ�/7�7b]���=�~�RMxқi�^r`���v{,�j�j2"V-�g�8`�����)J�)�
�1t1��{�X�k�ƞB`�\�+G�+��k�|~_�^k��e�&�̍1��_%&ZYʺ~F"�T�GN��ɬ�k7�p�|+�%1�����-�5ds>_�vY�ڮ�bsl� A���ϣ\f�z�`Q������}4db��]9r>�s�n��Yf���?��Y�ecr"�e�-o9W�ڑ	Wz3g���R���pi�馗{�n3r2���+t�V�B����%`zA<$\��k����p��&�S�ujĜRWE��T��se/n�� �x�k�T���0��&ZYVi`iQ���	O��]��i6b�T�6'
�84F��C[o~/���ed�7vv6Ic��R_<p� 8r2IVA��/ l�|[ڋp5�|�Dĺ,��{��C�����f���7��E'D���	�, f�~�᲌W晗�7�8��L^#4b�������W�?2U�7�Y����dj�F ���.E�[X7"f�,�*��T́d�;�$Lo��\�r*��5cs�/m81e��k�f�Z���Z��I��r^6<�Tx\p�um�m1�h9u��BU�{B�zʹxf�eK��Ͳh��l�@0��&��<_lN���:8K~��� ���z����4p�qs_�ۿ(1�a����uש�b���B�����Ͳ;������"6s�s���Jd��3���)���L�P�$�-35�2��h��c�uQ�9��6f����z/0j�Ĕmz���� ��u�u��M��p���n�]F�Y�����Ōf�,�fcc���Y��@G�h5+��l�65��?�O�$�7�ѥ���ɨ��ݪ�f��IZ��8�VB�6%��:`���������p�oy�b���|�XaE���b�9�$��x>+h0n�ug�����L��"���ʽ�WΚC+�,[�5:��
�Kc���>����u��Z!�����+0I��7n�Ț>bN�ͣ�Ā��*�����`6�G��]Mf�@�r� �,��9D���g�9Ћ�:P�PA��	�, ��z�Y	0b��́���>�g	�Y�h�9 b��5��q�@>�:L�����.��I�w	��Mב�@������LLݚ��*��55���[s1��$;oՀ�-}]��Y��osG@���� r��!����@g����Ȅ'�r���7�pB��dn83nN���G�rFm N��0~��j��bY�_��k/f���j���̐&�~ٮ��3��C�u�f��_��$q�96'��/n���'ѭ��&�{�����*���9W�(�s�G�+�w7r` �F���:�[�f	�j��G([�9�9('��j�x�]i1Iy��
?��,�J���܅v�Q����s���Yg5p���A3\\�����d3b"�e�n����X���ͅ�j�T��řg(��kV3�X�6^���Xg5�);��:So��$A��m�g`� �&I���Y�`�\��;v��Y��\�1�-1b�8u$�t����p�7�t���(���3b��q��gY���͡[OfM��Ҹ�0� ���p���R,l��arg��6B���f�*�Y�� s U����RKgi߼X�����*Nĺ���Ey @ӥaJOF�z_Y9$���l��lZ�gm����V}d�X�n����nY/dܽ2�M2���б���&�zN�fV<οSx����T�&b]�&ټ���C�������A����I'D��%�_�0��B��?���?�:_�E���%����l ��X̙�nn�%#��W�5_4�p�6oj`j��<�*L�c0�>I���m����p�]���f�9}��]w`8B�[^p�'ө�f���@�A�ʭ����Ӌ�"G�F��x42պs�|{61d�Uw�9�/�'E�_ĺ}2p6&G�ذIX���l�Cs!��P?��Í�N�:�&{���|�bΊ�m}��o�	O�_����<^2�
:��8�)h�3[�KM�~��(������[0��n�8�c�[77���-5���� ���뎮#zӛ �&�_�:2�sd�_��̠��j�9��}4l��Y���1�oB�69d�OבY�붐��eC���ͅ�`��d87cf!Z�m���$_f�\�3v�j݊.�.�ݤ�wx�W��
�L[�t��jذ9�u�ÉyQĠi�՜���u81�ǃ�*���m�dL֭�	|��߮[��Kxc+-�LR�k���2���cf���pM���nf�pG�D�����z�9 �Y�I�J/Z94�p���:���V6I�#�]�6nذIr,R�fVj�!�,���e����X2�7ux����饺��6�����ˆ�9�A�|�r6aJ�f!y�_8-;�܂$G81�Ѕ��F���5�y��Q���4,z�}�-�e�&�Db^rڋ�Mĺ��̕ZX��܈	S����2���w۪#����܎aE�[>+�kC���Q��G��F�����Ь2�1;ul��d����_�4�R�~���qx��F8�t�V���Jh�\���"N�@mJ*H�<a�d@���F�@������=����� 35�g�^�n� �sT,�%�9ke&a+������r���+̨99�Āۺ���܀��7�e�a9���f�$Y�f9�a�Zq�z�K��eu��I���7��:]�Heŧ�"�g&7d���Q5�s`RS�43�-��e�4R;9�s�n~i��oF��Nw]�lw)�|م��6f�Y߫�
d�1c�0rEW�1�L�fM��ecs�t�{�l~|w�,Ss���vn�c��̧���N݅CMXR_W6�60��9������a)s!��Bf�Jc|�j��X�G~�(3l��6.�l��/s[6��`4'��h�.��|�q��Vb��1S��!ΓG�#&RU��t�_�kxΆ!-�S{��M���ss{ٰ��rb���#{�Y���erN;6r6��j���P����tؔ�$�b�Υ���� �ĸ{��Wr�p5�4l����9��9�c`�@�f~2K.ZY����9g�0�����9�ASQ+F�b�'3�ŸkfY�i�QS�^�u:�wϜeu!�+Y��Yjb�)���k��/�r�wR�sw��v��4�����!GM������g�&RU�z�!��������]�es6�9�wI̡䪐��29�������C|��`%�}j�$/���R>��T�\̅��9�Ϧ�4rМ�h��eQ�̠�Ɗ!��Q��Y0g���.�E{E���� T�~y�$�"�L]_.K�j��rU�VK���s�.�Ӓ�F�x35�f�_�νA�x�zg�ꭱ�l��������
�	�����9U7db���^���
O���A�S/�ç�a2ɲM�;6���ԛ��iw�tYk�;Cج47]�H؜�8qeK�0��7��f�����9d�]�t8_{8�y�a#�J7�:K�"�[���`��:�Y S"�m�f=�71nФ���=]����j�� �;zt���d�U>���/s���S��Hj���nxȎT�rӌ4\72+����Hˆ��O9�:7�)0��\�+{��g��m�͗�W��v�,��Pd�򁘓aM��y"&iؠ��Pc��a�2-�!���	+��ޞʹO�u��V/�Gq�VawQ�Ɣ�wn��!#���9���L���I���\j51�^�w��a$ZY�ge�l携؄%�!�p�ᥦ���:�ȠI�_��FW}bN�$���{A6��+�l�$���:�1#��(�������ec����#(5��R`[_3n�{Ĳ�z��}9˲�d��+h�<@����M�z���nf<���Y�3D�ʲa�F�qf� ��,p�ԛ_�UX��^��i`6��L��qBj;P�PA��	�, f1}����,�B�j/�'.=C�-�uk����m�+x�Q����g�}8k�&c�uC�f@�6�Yh�-�����lej�D�lj{9zx�М�ۯ����$��B� I���s���n8]'��Ć�aA��]G����M���df8��M\��s��9����XW�;t���|����f
��,E6�|]V82f�9K2pF��
�%��YM����]3�G���K2�A�x<E�^w�"ǆ�3i��YX�9h��h���υH�A�ԭ+����a�܋X�rl�"�m0l�p皱��8x^8ذ� :X2#f���Yu�O��u�[>j^{�ΣV��9y��$�_�#���QS����萵��$�[/8s�nLL˿�'��21_�r�i�#��%9{ǔ�8���	ɠ9Xm��] �m�;61»hnѝ�Z�	���U:=�E�&<�O�\�l��i�m~�b���s����͹���dҿu[ݖ��\H���o�\`3�Y��uYbd.^��l�X��x
7j"֥�u��X�a�.�_B�y!t��������	3M�[�6f��J���9�!0�6�֩F�F�y�6�h9��r��I�_�p�܂��k15���Y�kwn��u�8!�(A� ��I3w�0\����bY�+�Ԁ�{ਹ�jodkQ�t�,g1r�o���S�Z�� p.E�s3�]��;O�pr��n����:8g�u<���D݆V�znj�fĈ�XW��m������I氶��!�L�m�ը9�!#'���*�0b*k�b��&�nY�Y�Ǹ}��t:���$5�v1+��PӸ<��ͲcF���*7\��a�Z�р�H��������#�m�Bi��*��VuAu�����wa#s�ɰ�:4��5Wsp������Q�ݑ�.�{�od�'sIа	O�#�̀71Ѯ;������bK�]��^p���]vv���<� �{�,�3f�f��C�Z�&p�Jr*
��<��o���yIj��tÆMA�*_�ͯ=��o�e�aAY�p�ȹ�I:�04C40�z��:0p^q�lNL�#�:Y�ȉX��d���v�Q��b���M�S�e�[9n��I>��GN���o,�9�N�0�
Oݶ�1I��V�p?J�L��cnR����b�����pC����j%��8������uY�������5��8u �5��q��qBj;P�PA��	�, f���9��cf�,�n�+�{�j��h��Z԰l`����vw�pi���d�&��pqj�,��U�&D��|^��}9l�$�5bV̺��#FN�����:�y�#�l�B�ܮd��.�����ۦl�|n�MR��o��mw;6կC��c�QSv 5#fc�cu�D++>�9�-��D��	K��n�1�SF�|b���n&I�Hub��lܘIBm��{t��A3xB�L�~��]]w��'<8I��|`6,��*0n�߱x.�IZ��kp�Q�6rਉX�r�^%5 aJ��u['8l�u�ڳY�nܠ�n�g��[�G̫̘1���^�j�F#�F.X3��y�u�����K=i<6����!HM���v��Y�n�$�;��So5�T�/4dFQ8fb��`�펈.[�e�� ��������6]w����1�fb�v�x`�HԺL�E%f�N�mѨ	O��Y 7���>5���q)�{����9^�M�|I���-�+����d�I����%$��@[E��Z��M��w��l�FMĺ.������KP�RZW0gU-;OW�L&�ԠY�uY�S�M�^�Ħ6��MR�S�-'�iΦ�r���r�&�~����[-�˭�?��F�o4�N'D��%�_�0�z�z���Ŭ��@�\ݘ��������m�����p+�t��y��e�7j�$\�R��3�� F܋i�p�NEj���ɬC���1lذ�j����s�m��#��^�`�)��e��N�I�sw��Īp�	5l�x]�	���]�k� ?���[�+��_X�73�����9�t�p�P�/I��?��Z81Ts��z���&:�0Ќ��c�²n�=I��@�p9qըQc��2&�&��&�����felή��a@LJg�1#��Kْ�smց�;eb6?��+��,�ћSv��o����&b����h�N����2�ls`6t��a�ܣ��Ь̺^h�M��$��BO�ltA��X0K���V�4�)[��%�`\d3I"��Y��Nn���4���f�rQ^v|��k��`�xF�@/9rk�0�*+d��\�r���nd�,�c�8j���\ݼ��z���^Nn�#�ys����65I����J̋���*��2c����_z���)[Ж��3#���ރ��!FM�un��÷���TZ1#�r�\�r��21eb��y�펔)S�Λ�Y�q{22h��L�v��
��BM&F�+��v���e�����g�hԄ%����� nܽ߷{m��\Q�N����x�$�F([����h�Đ΍z/���)c��&�Ͳ�5���X�u>�����z���a�,�6s�Ĭ�%S��[�st#1,9ܯ�J�$����k�-5p�$�?��:�TͰ��ь���+�$ssE���N�.+t�3�L'D��%�_�0�b�� �e%Ĝ��rqs�>�8���V���kU�L�.G�M9ح�4C�E����1&'Fi3k�d��y�BɄ��$�a#����Of6pJI���A`nn��J;8g�
^��T|S�u�=+�\Qs�X�;�2n>-�n������>�l�ʷ%����l��e�|@cy�	O�cm���U�Lҧel�ƺlJ�9�L}w7��5p���������pr<���X�}Z�jĈs�����Oyp�FnĴ�+|��,�%W4�F�g����^<S�f����ųBΓ.��5Qv8�^�k7e���-�$4/4��9|<͏��l��&���-X]8-��Z��۲�G�k�WJ�!ML���n�}�pw؄%�a����\�S}:��l��a���WE��k��m�%�)�K�)[������l��Ѫփ�Q��W������	���uF3�>�ԗ1�2�O\2o[^�3�!�UJ,���@����1�u#q�X6�g�Ajف��sxR�j>� s>�1�k7���C�*���>��j�lh�t�"�)��v�����&Y@Vty�f!s`6sj/�+�,sϽ>�ܔmͬńE���ls;����Y�M,�̰\�J���Q1��y#Yh�-���6���Kau�f��[�L����G��z�n:�
�s�����oi�,DO��N�?d�x׉)u�R���P�����Yǫ'����ZX�吉XW��Es�13@ '<���z�� ��?o�s�-������sr�1Cf�N
/J��c�N�\2=��`�
���z�2���2]��_�dh��#U��,�U���?S��-��oR��N���u)���mIG�+�ѐ��&�,��i�~���9��ej�	�\9h�eG��U7`Rp|��Օ3�kՖѲ_�r����pVaO���*�0��
���e�u�;����G�C�^L��3dCgš���}��'��q��\nf�̡i�ǿɺ�t$>т�&j]����[9�5�I�
�ە>��4���7�K8��Q�ܬ�*�O!2I�E�cF�a�2٘��Ϫ�C΁�rna�s_��&�x3'���,8h"�e�/��f�#j]N�������
>�؜�j��)��,۳u��T���t��A�ToU����o��uk�Fg�(&��Y��ﳙj�z�Q�V��uwS�qBj;P�PA��	�, �b`��Y�5X#4'��N�YF`n��et�� 1SÞ�rn�1%�����W���;�g�W3���]����/�Nڻ��s����ή;ظasҳ9�$�3H��E�f�����0dRy�p�s`�3�o_�P���n��d"ו�]y2�� N��qs�D�	S�@���-L���z��t0O�:6��M���FN��u]���w�I�-�ͪ9���.;��L>��o�X�us�*3c�az�1���R]$Ƒ�u[mt�ʟ9�"2dN��&G���D3áČ����[�C��
����z�9wb�R�`�����M��Ό���u��1֝�K�;����>J�i"��К�W��-7�!�0`�b�u��9ĩ�FL�:0�ո9@��nи	G��݁E��\�Z�����y��
F4������9А9�ԠI֭�I����m�3�Y���s?�ρ�_0'����Sw�.�!��Z���;��KVMR�u�Cf��F�Z����B��]lb�gs`_����.��qgȹЈ��K��[8��l6�~[]Q5�9Lu���^I����q�f#dV��&R����!��R'fى�+��Dܚ�Y�˿vf�D,˾���>؜�n�|#f�^
�%jj�3mse7�Z�:0jT	k_��9 ljA[��-�Cゾ13�Va�����JBۛ�7~t��X��/���G#�==����l�E㦭�|hj��a#�(uf4�zi���Q��[̉���hH7�w�\�h�n�×��SN�op��
�Y�E�&ZY*���f�
�	Cꁞ�Iq�ȩ.����s�"N�@mJ*H�<a�d���s���+#�Xz�,����/��L| _�l����Y��s�1f�1tb���Ժm@�z�	���e��7�(�G��nf����.LulVy�>1`����pf�_פo�}����`�ep��ˡ&	N/{��޹K�L�eF�:�ٜ���,[��t(���d���vW�zگ����s��Ɉ�Q{���]5��?���$A3Rٝ�J]�d�M�9��7`Z�e{fm�����dݺ���Se���%�����Kq),�u���D�K9q޳��2]��u%�ҿP�k˺
i���,,�$�x�N��#z�F��>�ށ�g��[K��dN�N56�f�~�&����plظ���Ⲽ6)i��Y>p����nǲ9�VJN��7�8n��6����� ��_�쿗�������Y��<�0#���J�1h"�e��ez�Ɍ+�I�27lY�9�p1w}��7��Q����f�GMAQ��<�&7��jb���B4�N��B2ɗ�S������f�̠�X��_���J��Z�ӳ�����qS�h	��ɹ�M��s�����M����Yh�<�Bn&�޲[f�B8�ܙj��[˅h���L���A��v׺$��Sv��e�8!�(A� ��I�aB`��9�~嫾d��#lɢY���ef��2��ȻP76Z�I��p�ӃϢ�B�N�194��jr]�Ԙ��t8�/�D�b�����j!R����]���[ʨׁqs��ͩGM��E48��[�j�,�e���"�[$&rQt+b��yٌՇ�w���3�>�^=qbݡE��b]�3���~n�����Z�b�,{1I�Á��a��	�26��3�搼m���Y�j�ߍ�Mx�6Nf]6�H/�)[��$g1������FHnن���z��
ٖL�e�yp2n.ͪ�i�&��vbb�������}�&�����j�b�.��Kj1�a=���6�l=Ǻ-@n���-��X���11�Ǘ���+ ��4��7}�Y��fT8Y��e��0j&Y�i7'��E)��[M4��z�Yr��mv��jޮ&ZY��.�KeYo<bYI�F̝s��F�-��f�c8�25j�����-Y%2=7�:'��,�_w2��fR�"7�n��2I#��"Rs�$�|{l����fi�!��d��i��M�t��HΆ�l(��a��gf���rΒ5�"N���l�lp8�hαp6�&���ê>�M����"X�7��&,�W�Fl�|x���|Ѕ�f��Q#���{ov�I�"J��A3�҄�&Ƹ�v�.78p���zG߰l����G��!C��heٸK�h�؈e95���2+��M���-XC�}��e�Jb��4گ�&�^�g?���]�hΎcB̈��
�Wd�$S�~b�t;9�SK=��Z��"Pہ�
�/O�d9����������[d��#�`-f�mdkQ��pG�;֡�8{�XVjV6f�d7�pY�j�<��ds��26'�9'���$ �����#GLx�ĜT����N�lϕ�139>�Y`Ρ�vCf�X��&�*2]%�T=�9�צ˞̝[���蕹�lԠ�V�����~h�V����;ß%~�H�{�6,�Ii�l�,69�}���S|٩F�;��I@�ˆT��ꓩ`zt�9�o�3I#��_0݈A3���qf9/�CV��~<��%G��he)W7��C��'�_��ef�ܟ��5�z�7���$�Vf��0dF�`���U��
>>���������3��23OxHX�w��ڻ�r�l�P��b��Qs7We�[���Ⱥ��ĕ]���f3^<9g�Zn'��W�&�[.S��,�K���E�؏���~������QC��%�MxR�97�8p�|l���꧿��G([�V���{)�,�Vd����0/��6.��:�ϥ);[���4�X�oTYy4l��������@�3n��9�՜9p�\���݌��u�>ō���j�iگ��nb��dR͇��F��`z��f��1s��I���75�~X3����2�w1-�Z��"Pہ�
�/O�dY�����sF5,�%��1��i,�C�Z԰�j��� �3�3�x��Y�uH���lT_Dg9��(;Ι��ɟD�}��Ma#f�Ą�l����0�[�fR/�dƟ�0��n�ٹ�ə�d�*�9��I����n�\���1�L��wC+W����0�-5�ʲ��p]���2_2aI}v.(j\�z�&����b�$�'R��Ά�&��mJ��l�?�oñ�L��~=���K֏�3r���I<�9h�CO��Z�O����LR�e����8>���V���A�-��e%5�|�OQ7��)[�k�f�?o*Y��/��<D��V�.��&Q���,�{�WE��6��~��V�,;����]{8-�A|N8`�$���pN29�~�yսYa`�Yw6qU�ơe�-H#�V7�����rsl������X���5?"�$�0s>��Wo˲�+`e�����^�!-��2���ߘ�u����|��Yҧe�`cf�3f�\��h��$<� i�T�+k���B��`�,��jn���=���#������d�}񟎇���r�h��qK7M��as���`���3 tc��a3� f�y�?3��{����S���l�B�`ؔ2E���� T�~y�$k�� �.��xZ|���=��gU���^�m63��Cۙz�Z��Vf��7�M��u��fi,��r;ƕe�9@�Ȱ�)�>����ө�`e�M��e+�0�񃳚a�cn��E`R�����J��D++����tݗ��Ð�eG�Bof�gT[��!sp;�%!�5@s�Y6�����m�o�&�dʖ���{l�K��z�ĸKfU��h�S�f��Q�c��I�e�d�f����r�>-���mWNJ�]�1��L��̯E���A�h�����3Z+b7<�xK`�.������'Ǻ�HJ��l��z,�cFM2�Y^�k���!����[�I�t�zL���la7��`ܬ��3)��A����R֜W�O͋gQSߖU97��p�;�,�p��$ɸ�W��Zv۸{2llSrJ�RF�p�fi�Y��I?B�3�]����_�c��$�{٪��)���ƪ�9h-
9l��ejܫ��A�L�R����F�T$�98/<K`��I��25l6�f]�r:y���b��rY���9��.0l*��Wō�X��U�ڹz^��#��
g3�;�J{9M�uFc&��K{%V��&'bY�|�NB6�V���$>�7��4hƑY�.�X`�ZG)[�E��iבL�?�N�a���N��{d.��ի�Z0OKfL��rn�a�\�heYd1�s)�L3#'�#�G��Ɇf�)�W�	��@	B�'L��ܧz�Y��v�p�f�-�8��S�͉��Ϲ�nfB��r��,���dd�������?�.��f��uq�κ��p�ș���ϳ���M�l�<�2X���A�u9�9���.jRq^�f�,t�ͭ_�:����Z��f���n�;8S��O����d�c^����A4ZYqW�¿�޳|��	K�v=/�#b�д��3f�Y��$�٩v��!cN�p�_��ey�����P���M��(erΆ���m�$R_q2��(ږ�q�|��C�l���,�S�he�'4'��e�rX$aI}��9�-�C��)#s b�����N��댽<��fXs�C�*��&�x�n~�.HG�{!��Z�Ϥ��c~�-��9�z=�,��Y�ŏ�ƕs�$�"4��o���ɡ�d�5�l'��UӢov�����wܬ��_���8�U8��9��r�#��g�*̰�|Zf���nF���V7��͍���4�xٳY�Y�����x�� 91�#����,;6�)��6�.d䜄�ajN�uws.��bn�e��bb��n�7��w�,���^HN�%�NxR/W5�t����23f�j2�f�M)S�	��@	B�'L��mY����/�{�^4���,,�sq�Y`Ο�8�&��ҽs�\9Cϲ��B�&��e+�����-�$q�����1p��sd)hf�LL);�%�A�(~����`l�Rį+�UZ�j
ې3ebFٕ\����UF�暮��=�n��e��/�s,���{�/)2�k%g1-`�_���S\�֕M���b�o����ZᛸOC�a��Φ���Oi4�l�`u���D�3 'f����(���<�Q�0/��i3OK&S��F�u<��Tԭ�ldC+/'&���XA�:��i�Z��f�=�^��j�e�%���w��}91>�9��v#�2\�5:Ly1���Z��v7f����k��d�l�&�L"s�M����x_�r�,[�����ELU����]����sv��:;[���i9ұI�>�9-N[0d�� 0�#FL��u]�y�ٵn���ԟ���=ńDY�
b�P��ź��o21*����:�����	-�R.?9h��e��o�NV����v�W#'e��n޲�Zhv�t��-����n�����p#�ͺ/0C�U~8�<-b|�P�f|_����\Q����I��*�M��g#�\Ќ��IL��� F����Y�E
&bYt�D+S�	��@	B�'L����fy]3č4�N�Y�er�·��'X�v4d��Cছ�r����m٥�E�:��y����Q� ��EΆ����ض
��ہIV]hg��3�8�TU�X���= �q���{r�9Wֶ��������I��l��@���m `��U]���;�v��9&Ȭ'��@�I�f9�A�4��w��f#3e�d9K�Ь~��b�;9j�MM_V�����Fb5dЄ%��.G2d�NC��f�و��1��g���f��{�p3�)i�T/�g"3��fЬ���7���lg�I���n2C;8��86�$����I��f�����Ԉe�'6`����'s�Ò��9��Y94�xݟ�['9h�Rv���{�%M�>�s�Q�&Ɗ�bf��.�
8f��L�$�u�b#gck�m`��l��:�9�Ȅ'u�.񍙹�`�d�(��v�����&Y�63��������]�ܘ9��Ԟ	7�]i4Ow�հg�B�����`i���|������s��9��A��۴�ie�4[�n��C�{�&Y&���r��#'�7*g��R��e���1�겧>�Y0�,���D�-Xo2c!9�21�8�]x氤&#�0y]Wc����L?���|4f��S���#�&ZY$ʋ	1ʟ9
�6Z;6�u�Z�ef&���z�$�ū�&,epV��ވ��M8�zF�Y=7O��N���-�~E�s�rʏ%�i���ݍ^��Lޕ�:1���Q�M�su"qELZ�F�`�4���h��Z�!���$� s����+Yh�0Kw�����f6�Nk'N��Q�OM�1�Z�E%F�B-&< ���\?1�֡-,eK�e�g�j"rCL-S��nO����㠚�:����kf}F��Qs=�1�?Q�.g�$�I��h`C揚GO�
\G˺XVD(���v��|�O+`��%.G�����!����D�˥fAZ~�fR?��g�/�p�F����2k��<��?�$�fs�^��^爰&&2w��2#�����v�Z�b���q��ca���.�G=��!�f�,�h�ˈ�22��<�d�DL�ec#f������f�̬��K�S�7��&�5W�l��ج�鑤}|���9l�3`�$i�j���Г�X'��Afm�D�%so��5k�|+�F3��	9@[�r��^��e�ݸ���
�����Q�6� �F� A��9Cf � �`y �s��l&Yv��7�1�ڧu�ؠ�^4aI|�[97'�e��]�sh6�&`ܤ`����?�L��lU45��M�&w�<\��{]��Ԭ�wp����md�������);t�Ybw�ɲ�Z��������I2+�rG8��p����!��.�[�C����9��,q1ɪx�/�lF���ݐ���f�Oj�k����Z�y����e��UCsБ#G��$�7O�
��ӡAZ����b��Sw��'���d@�-+>��WbF�ko&<��l����:����~���u��&,en.�w4�%Mҧel�͟\dԠ��i.m9��8ͧ�̰p8ؑI�oA3sh[��i##�e��ŪfARs�:
��8�+s��d\)��v�����&Y@nS=�p3�6�f���cN�s��ç���o��a����mލ���9 &a�F�딀3B_Rp�n��qI���n�$���}�"#�u7溑�fR�}݁f���X[6]���d٣YjR@~��qxٲy25���L+��l�L�����M�l6b�T㏝�\�'i��n�9Q����_2�I�N&1�4��`��u9�/��I��1��9��tz0��F����4��=�_`�t�N7l���I�4B; ���=������i�~�$,�뾒�\�j�Z���Qs�O��N��C��.����$}�R�Ͳ_zG��:����f����3u�e1���gL���뺯˒��]���`�d���h��=7s  �.e�ɮ��>���_Rj��73M��<�և�{����l��W[N���C���RM�n�Vq��f�%܏R��nN�1l����R{fР�nY�܅�np�dW��j�2r��e�,dn�Q2aJ��������<����)g`;���sb��ʬf�����N�M��9kω�+M!�3Y�N,���،�r�.���n^6T�R�)߁��&�ʋJ��~,.8�j+��䗳i1d̄)�z�I6kU�Sgt]�nnq�����,F8�4ƿu��X��J���Lof��t3_�m��.�ep���_�`��n�a�&b]�ﲭ�B~��1��Q����985�@�N'D��%�_�0�b��0��i�b��9,�9A�䞅�2As�"���۲`���l�Kϻ�h~�)�F,ss�\'5dܼ�M��u�ʺs$� :R�lat9���Mt�{�j�y̼JLD(/�|o�oQS�Al���Һ�s�X�Qg�Ĩ�����7Gn�n�`�q9�]�m�r\h�,�c�M���������,����D>��[h��Q�T�ܕv3٧ns�8���b$�G�{ 7K�̦��1�Ir,��`]��1?�1s�]���
~h��@GfsrФP�|�cfeR��*b]���{��+��Ƅ'����o���uK@�
Zg6� YgF��5g����5�U�x	'I��Ws}��ua2��r�Ir.Z��:�97#g�8['��9��T�!d�֕0�8��_�������I
o3�Cs�.Ӣ���>��IR��[�ۣY���ua��ef),�0�L��1gQU�O�usx3�&��;~���J�6�mf���ty��n��=�7I�#ԹY��܆�]���� &Gι{��3��F��`������V��m��ff�����!7π�x
����"Pہ�
�/O�dD��v�Z�YɃ�9�rϊ.��-�d6� f����S�M���Q�fI�y�b�+�g`l������}y,R8j�e��n�np�g�43b�e�r&e�ifܫ�c3e'�`���u�Ԍsˑ�Jm�*��~�n�GsĪ%�x��!3xh��ܰM��$�UCf�w ��.�9��E�f�I�O�����������K3���� 4G9����ξ�xcs ?'N�N��f.�PM��uy�9��r�E++>�Ws�����%���+����eks�=�UJ���܊��O&�S��u=���Ͱ�a�{�FpZ��#��N��&O��)i$��X��^�m�L���v5�����Y0�ˈL���%������f���D7c���~^��>���_�h��y�U��κ��*o8�a�21�V��S�
&I�ed��]^�� �M�͍��9�fy�R^ 17Úګ9�Ϙ�79��2�V����A�L�R��f،/h��)�k���2ɪ���U\M1���Ѓ��.�`��s�.�A��rs���r�ȉ�flٺ��l�vmc��ͫ�Ʒ�i��x�������٠�����V��_�x��T2fz=����xanf0�j�*5h�4Ck81�D(�s^,�e����l��� ��:ܬክH��jRpΏ�D�,�t�W�
Ò:
���2w�m�N�)��v�����&Y������h�̩JN�Y��,�vY�i�v1qiz]������Rv��iP�$7-�Rv,,��5v�&ʮ��e�F��ƌ��S��<:�uS�^WX��S��~����}YM7S��
�$Y�`b��,_2l.��ӂ]/8W좑�֩?��o]�kc&e�	g#k`�.܊��hn�y�C9	VU�I�{���/Xk�ƛc�q�Γנ9eѰ�̟(�Gj�g��Wl��p+�H\�u�����F���<��⮝+S�FL��fRŧL�%�-355�헣8WNjĺ�9d���ڠ��m7�f �RQ��{������Y��u�75W��ml��5<�՜�r������`1�R4f�F����=�����b!���71�Z7�@�]��=���p#�O�_2pF�_�N��6cfp�F�����f��u��%
fḀ�$�Ь�ʯ�&�c&b]滙u;ۖ�Q���7���>���-9`��5Wc&�~��u[1��caK��MnnWR��6\��lʎ�G����Q��6֟��M׽����9Nv3?�^�l"�e~������l����.Dj�^+|M������%�za;h���v��<;���u��(ul���1h���R�t��Y&dNZ8bb�-ͺ�)�+t��;��o��9��[54n"�ej?�A ͱ��Lx�+f����M��Z�Qcfa9�ĸ~���-b���ȩ`t�-h�z\��D�.���d%SH�4W�4�h4E�{�W�̡WL�p3r�B��!S�}��h��K�5[���l"�e��e|5s�G#&<�We9�A3 ������Y��=��E���n/<�/��N837~w��$�?VF(�;N��ũ}����(��|�C&b]�	�@`fE�	S��?6Mbܘ9���u�8!�(A� ��I��Xۥ�ַe9��� ��g�]�蕾�f֢���_�+SA�[��h�Z�b������������~��P�܎擘�u�#3�%�hp��/�*�x���M�,9?v1f����3���yy-�m7��"7Ȱ9͗�&А�����fu��5��jSwe�[5kz��T���sؐI��n�l}���L?(Cf�(��]'7�-�77d���ʅ�LĲ��R]/4n���	Or2���\�f�TYB���|�&Yw>�G���:3�Z�6k��L������"v���ڨ�$n~i/+3'�RS�^߃��\Al���Y7�pY�6M�͜Mg��B&�3d���>7O��[�痚�gGݥ��(>Q�������3���p�ͨ)���y���A�5ɺ�~��!�f����ލ��k�:5��y��9	�#�-]4j�,J5W/ɩ�uTc�@L�­�3`�O�3���-b3����.\-y��;�K�� ��kN&K��/L4dr�iv�쮬��z��||�Cu������$�[�r���s���)��v�����&Y@м�����`&7��r?r���Ɩ��� 3�nظ���᦭p3\�Z�k~<,hr������y���͔�qsW�j�qSvJ7b�&^nl��[�I��޳p>�섆sZ���`����A���������;��6k��]*r�;׽�]���JoJ��v�l�m��^S9�E�%��5p��r^v]N��Z����O��Afʞ��-�(	��z�\m7#�)��j�N�ùj x�۬!0f"Ue���Y���hU%�q���Y�[�[@���0j�.F({�V��i� �l�~eŐø���y)�.r��aca<��I��f�?��)����l@)F3����f}�D��|p������H��iWnR�O�Y�̭�FN�<��h���]�݌q����gEҸe��ApnZ��edȬ�Ž�f��`p���ZBd�.6�f�m��I����u�>n"Ue?��:]�lk&i��lY\V6�!3�s�_Ar��$m���mf��d�A�Hf3p�b~�K6��Yp���%S��3̺��f��%s.��G8I���Y72d�2+��ۚ]g5nbi�� �pn�heY����9h���7��B>`��F��g��{��C��ꠉ�)B���L�vh�F�#�y~��Lo_ �2qF�Y��Ċ��heY�q��s�.���/8�����.U�	��@	B�'L����b� ��`Ā����P|���U[F[�dn�	VÒ9�,���`�[odִ-6W�88��4�Y��l�J`�$�֜��uax@5S�����SM���X�58��Ͱ Z��C暞��B&�y��e��LXҾh=�&FLuoE䬰Y�q�*2����fa#'�G|�j��l~�##����ܱ��Su�h�mn�$��WG�"�3�����G;.<l���94��&�ۛ23lN8f�Ʌ�L=�,��l5�Ճ=�#�6�z��Y�+�ίn��nmj���h����ȬԔ���+�V'C�����f�n+'F�e�9����8K������3h�d��Y����������v#hV��x��@�� =��$t��rw󼇦6Z��_HV�/����3�y��v�R��u/��	go�K>es�9�m�$����8�S��s_{2}�kJ&��X0^ճ}�6�P�IB 1ρhғi�GG5��2s�TA�)x}����¹_���uZ�1��kp�?C��������s#'<�o8�,g�p�4#����fs�Ÿ��G�ԲIr9J�9���9I�_�bN��]��e�r�sb\1�m��N�������0͊0�=���v�,�qq=V���=C��晸y3n�,�`:���YW7:4`�,x��ڒX�%���@.���g9�>���V�S�6�63�2<i���좩A3,�C����f0�21wja:$m$	�Qʖ��LͲ=�bh��d�-�k1eOg��d��pq1܎0d���r]*0ی��I}�Y��w�ظiw�,n1��%ꦨ��"Pہ�
�/O�d��� s(^H�,d��E�CNf�nl��X�	Kf�wf�e��٠��]�+jf#��� ��n��{�Kk�l`u�t��-�jR�N��-���a1]��l�49�٘u_�l���[g3'������A)������
M����b8�7� �>�I��Z�_n�Z�8o�
�]��/r1��E�Q1���,�+C�Ĥ_s3��ͪ��6���X��>���뵆����Z[�4W00G��NA�ud�<�jmN-6���y�*ap��D��|=k�\�{l&L�����ae�JlF�M�Y�7�t;B�
[���I���-tb�bb�jF�!�¶�����4��A'��A�ݕ�E�f΁�=�ɻ��:{ɌM��R��9���c�Lxҫ9�Y��zP����f��IY���K���1�h8���ZM
��،/n6	怑�f������+砄&��By�q�M��s�c�R�XL/(rZ���u��pn63!2�J�^Wh����5_�h��J�r����7��e��pw�Ԑ��0���Bv�6SH�f%������H��eo���3r�$�^�p*G��J������&��rЈ9�/.7��~�۱4f~!;f���,�տ���cf/Q�䬋2�x�S��-J݂��&s���&��u}�s�VҐY0��e��������5�,��u24����u;6�F΂Ȧ�C'D��%�_�0��4�ȁ���`�x��"'�����F̱�튛����&7p	��6�M.�[7x{���\�uxy���x5�n�P����_T�e#lh��,tbB���a{��ͦ��H{�r_0`�\`̄H]T�#���e{8%�f�l�&	NQԉ����VE�[��$gs�&�y��������&z�(�G#&䈿�p�6O������<��C�}�(�Erp_c7S&�p��le�$���Y����b�lil�զ�1P!�����p��)Ss�WA͊�#&���Y��W��V����ޗT����Rp�
/7Ӗ�Y8����Ny=7�f�L���
h��o�Lg���}c�y�*�Y��ĸ�^K�\�k3e[,�G^�r��I�&�湗0p��<r�АY#3r�$�6�ox��,��셣fi�̄'�	Ȇ�E=sG��n���%KM�����Q� f�p1f�D�3^���/���4�z�rd���:-2h6�&鋙ɹ��&��S��l��%�'���c�mz��D+K�]/���LXR�9��Y�e�l�lw/7K�$ɤ�п��c��g��sU87�L	�6���hQCFM��ʖ�x��GG��wCf�u7�3��j_!7�$�9���� 'ZY���=V*d����*��b�����Ľ��9�t�P3@~�W|-����!���$`�aĸY��/�Lӱ`�c`7Bك�A���Q+i�I��'��J�E���73�4����5��M�������3om̄%��M���dĨi�]�ǒ�#JL��Q����Yh��1��)J�ҹ�`.�3nb _��"��7�\��k&Ƨ�ͦ�܆�5�,�·[e0�'�K�����8�W��Z��"Pہ�
�/O�d���a�0k�&`��`�kJN�9'���鶏U��9�ݬ�rm��� 3&��6��"��$�r��(���⁉�l�c΁lZ��);a�,�qUͤ~���f��E�,3Wq���æ��+��y�tY	̨�n��P1e�Ժ,���25k�n��Pn�D++>-��i	���2��=��_0G�Q>eg.�-�ȑs+�Rf����F�O��elfY��_��Iͦ�D��5�`|����LFM���'�0b�tٶl΢5���(0p�i�����V�rw��f]�~Ĳ�z9�Wn%����sj��321U'1���F/�v���a+x����,3�d��j]=9�X8+tٓ�@ɲUFsHY��O˶�x���j�V��#�f�v�.���f�ḉ!�]��,6�fp��d�4��<����T7<�.��/�H_��#�BzL �#�eb�Y��\�`�MxR7bݞ�6p�~9l߁�l��܀��s���k����r��?�v��9k.�fbɬ��f�����`��_96j������r�ĂQ�,�+f9���V9b����L����?������1l�h��dڑ��Xq.�qō����,�k`�p��Rۗ��,7�.`�qB�#R�<�B�	Țo�H�:j�$I�T�d
�|�u`J��a	�)�Gh�~nP�PA�n��=1.K��d�,95k�)9�X�S�����\o5�n�r(�8�T��geĚ��2�j昞',�#TF�?��Yf�3/[8';3b�DcO̩,��%��M���L5sl��ڬԙ~���J�4	Sa��E��[��͑�o&I��"���a,�VqR���f��ȁ#���f�ޛZ�����.6d�C3b����09f�6�M��4m#��Y�p�0+6l6�0���ӆ�0��ei��{ es����gzÖr����sCf��Vtcl�,��-'JI��a*�Xr�D̦�lv��	K����!mëY�ѐA�Z8�R����j/�':���GWR����&żn�j��R��caĒ1i=�D�;��mC�0�W�8)Űq�5l"I
gO�ھ[�C�.lV�ʪ�3�`�T�֓�F؀��l�D)��=\�K�p�}��M̢w���um��2|u��$N22jԄ�b�p#g�嬔4p�L�H4�P��;�.Ks1��5aJ[���i�Xf-#�`5�l,^�t��k�*[�Y96�85�3d�,O6dn۳c��Z.�0�$�ga�%��f����<6aJW�֨i�Y^Ͳ�Q�݃��ͺ�Q#Fͦ�p�s���3fܐY�Ų�nF�Q�͆����%���fk5`�5aI_���i�Y^����𯅳X��Y7[lu4��"�M%(dF��s9���BcFN��4u8+��,���rᬌn������č2bԌ(�m�� ��2f��E��Y)0jV�;7:{d��G��=.��߂��v�?�=X��N��"ԹY�p�,�x��݂.��a
ua�/Z��ʌ0k!ftZ��}�A�/�e����٠�H5qLWe��;|ZE��pVF�?r�pV�Y��B!7ֲu�!�F�46l�-���;��,31n�|�u9bn�6�P����&��k�e)�1#̒^�=8R�C���p3h��fV�G�IS��2z��=e W����GN��0k��b��ă;����1s�.���H����n�r�b�l�#F8#�D�"����,y8+ìe�<
N�͚���N1�A������*0Ԡـ�H5qd
We�8�Qs(���U��q��폜:��a�:'dԨ��o5�!G�4b֊LD���j�i�&��#',R��2zMT��Z���R��2�Z�I�14f.�H��ҫ�2r��pp�e�A�&&C��Df٪Y��&�a��^CfQ�q��Y��ȉ�X^M��n�,v7뾶p��#�zj��j�O�7hȄE°VF���oX+��Y�pV�Y�8i�,�u\�dR���e]�����_�EoF0?Ĭ�±���Y^�f΄��]�w��s�"��>��l�*\�,�(G��o��t��R.q�z�43NDWx(Tm{���YH�Ė���,*�?�O�5fVm5/�&��4p2P8[{�7��T᪌^��5�܍�E�(Մ+u\ed�#'cax5�#5j��46��DD���b-dhܐ	��a��^U�VF�?������ 2j�Ċb̣�1��h�ZT�bVT��&��YH��ac�p7�&�-���k��Ոq�pm��p����n��a���Y�(���q�f�Ԭ�y*F5`�~l�Z7b����6n�D���+\��k��M2��2��QS��2�Z��l]�#p35\���p�1�&<d{j5͢/��+��5uX+ìu�q��4bV=\d��	Üzq��&Ԅg�Q폞:��a�:gg�:��e-��YK0pV��[m
�&���̈�r�.��[H��R��ca�9\��ِ�(d
caD[Ð6����,*�'�6�af��\Lgz����)�mZ�j�YX�[N��8��T���K�D�p#�9mëY�АA�Z8�R�a�5�̆WtN|s+��$3+���bv�1l���i�X��4X����@�pF�5i�X^��\w9r��KGf5�,���b"�L4}��<&gyo�F��Hƺh�uc]D�� MëI�4dԬK4����7#�W�Ɍ�#&�M�e�"+��4j���Q>L��KؼDN��M�)qled���gex5����5��f��q�F�Z���w�V�:��43p�C�pF.��oX+#�]�pV�W�0�j1sY=5fθ�и�S�+9p�-2���[͑��QJR�X��xBɉa,�hk���,�fY�(���q��"�S��И��̍3��f�1�$��0F.a�1��j6�0��Qӆ�0�����z_�#	�'L��� b~��cӫ����-20pV��-�D��p��K�[
�p9�����[�mB���3'�Ux|��X_�LaU'�6^y0k*f�l
�
��A� �N����bZ9�j��ᬌZ���u��DaJ8+�������q9��D�؄p��>2f"�+֘�(Tӕ����P(��52�{�b6�,n6���ĳ^3북p"�ı>\�Qk�ר�J�pUF�=��X^M�
gI�q#FL4��@`5W�{��j�e��{��M��8��T��������q��m��6����,KE�8L��-8d��� �#�%qƇ�0r�������0F�5r�0�W�8|�Q�&V*2kw-z0h�F��*P8h�$(�%�͠�Z��r�0�(%i�0F.Y�i&��Y���i�X^��/�����y7k}����9�np��n�	�$a��ZU�0�E�-��a,�&q�a������m�˺�Q#G̊lL9f� �c Hͪ�Y!bF�.�	(��Bcf�޽^���L�h޳ݪp9ج�����o9j��#.�i���2p�(0+ 4��l64�u��^׺�`���@���B�����>2hР��W�f��[6j��A�&JI��0r������pnr�	Sڸ�ȶFN���jGF2j�<�0����T�v1+Ԭ�1nМd"�ukj�n�F��#'D�bE	�!P��+c`�PK���eu՘9o�B��
!�M��K��K�h�Ӎm JI��0F.1��5�B�y6l6�0��Qӆ�0��e
D�w�7�fe*,�ol��0��Y9`���fݣ�����%r^�&
,��0��Qӆ�0���A2���,��͊�Y4`��
Y���A�Zd5#��鿬Vdo��&RM�:���k��ٰ�(�get�#�ge������uQ٘Y�5Ss�Q�&h
��kW��Ֆ�0���H5qz��2z�ר�B�pVF�?r�pV�Y�8\�!���&V��p���E �Z�كS��	8hd$��͠�Z��'#�M��4u8+�����j"�1���폜:��a�:N�uT/5��_����bn2D�_���jCp��n�	���,�\U�pF�7�����qR����uA�:f���SP*��6�݈sĪA#��H5q�We��m��M0ket�#�ge�����5j���h��(9bܠ�fd"j�TR�N�7�9a#���k�j����G#��a�:|�w^�|�VA8�p��Y�� ӡ�z��WG���D��!A�*�׸Y�cE<��2����0�����~�7����˹�b�pcn�;���H5qz��2j�b$�1-l�mC�0�W�8�Ĭ�2d԰�$�F�V�Z�As^�Q�5h��9&�as.��&RM�a��^sz�����UF�?r�pV�Y�8Q�\� ��y�Y�Z��Q1rJ0r��q�:1p��	��a��^U��VF�=��a,���8g��nȈi�I��u�Rb�l|m���!f�̬���Y�f��e!7�R�^���E��}4��N��Wi��Vw%��7��D�k]6����n0{g`T�y��0����x?�W��n��F͂�f��fS�LM
��ш��Y��e��8�WeԚE��c뾈�6<��+�������q�53��v�0p�h1r"j1�����uaCF�8a�>��Qk�k�ʨ��A�pV�Y�X���3k)g��<	7[l�D`���ɀ�1\6fY��l���H5i�pVF�a���`ǩ��q��폜:��a�:�E��j]Va�<��M�٢/�S,]q9��9�-'JI�>a*�Xr�ȼFNr��2���H���j�4d6��p����S�H�lxE��T��Q�x)yȘ�4[��]vdİ�T��ge��E��r"�'���폜:��a�:N0�ҒY=0��(p��Ȁ!Qo1r��Y^[���&<���0rIT]�Y���҅�2�Z�I'��7/T3��2��:��#�1��#ǌ `~8��z+L��م3!�pY(̬Ի��9��o�{�[�e�fm���o�m��k�f1�Hs��͉�΂�B�L����ؠ����W�����lh����Z���f�����}�@[�~��[6j��A�&JI4��0b�m"�SDͦ����$�P��p�gex5�#32����T�j;hN}2ѴhXR��7�9�:��K X+#���Y^M�>s������}�f�حиpj #L�rs��,�5V�fc��&�%���k�lv�]��&ذ	W����GM��0k���"�7n�mm�T�X�k���ԍ3���6��$N�0F,ڽ�Lr��2��aH���j�1��^XqbfShجv��_2�=5�C����$�2��QS��2�Z�'ϵ횠	��k�C���F�5��U|et���ke���Ù1r�ȉ�9p���r��VO�pmn��$ȵ��z������F��T��ge�2wZNr��2���S��2�Z���I5@� Y�=0sl�f7�f��j���l���)�c���9��L��La�0�
�����¦�2�z����F�����f����ٔ.�o
L�Id�p�����.2�/JI�6���K�k=�D`F8#�9mëY��0p���&�:���ƌ�_Or^��s`( ^Lr���4rШ�R�w�
#�,�ͯ���а��/�hk҆�0���IGdV�4ٵ3H�DF1r����_r؄7a��Z�\a��l[d��0���I�q5ѤX{6rV
�b^�hdh�߰���#'xgaĒ�dgaD[À�0�W���Y.n��C�F9�f��Y�����</���aF�8h�,g2b���i�X�d㇂ue#f�0��+�lk�a,�fY�8yѬ�8� g1l/����t,�/�Z��ͺ�Yy3QJҴa,�\��b�d|#�9mëY�6$8`��kO̊��7j�j�l�F�4�)48����\�?�"��ᩋV���� �������E�-I�X^M⤺��g]��f�W�Lg?t��w��A�w��YG7b���P>\�Kn�&��a,�hk҆�0��E�����F���Q���r��U^�$x-��Q�f��i_G�0F,Y�`��9D �0F�5i�X^�B��pY�S��&��W�|Úr1.v3l؄���"���a,�&!T��r+ F�(�_�oڅf��I�0F�5i�X^��(I�p��م/LzǗ�E��������mC�0�W�8)Ŝ?n��q������Q��m��I��73O�,0fԨY�V�!-BM���2j.Ks	.�p؈�'<��+�������a7p��.���o��fc�?�^���Y6��L�����2j��bGN$��Y��0�ge������gp�'{b%��s���;�p���rS��rn�l�M�^|I)�T�d�j"�B�������Y�8Yo3r̀a�̚���5�}N�徇��I/&RM��V���n'�^ᬌjR��2�Z��3k��M4���[땕�>h:��W�$����Qs�l��<�&�|᪌^c���d:�2���S��2�ZǉBf�F���]���Yߚ�81���/Z�Ь�ei&RMI�V�f�,4��get�#�ge����z��b��~O̢"�A7j&�.�3L��z+�f�n�R-�$�a*�\r�E�cat{#'ge��3��'p���ؠ��fj"8`��hr*�A���9��FL�����2z��&�Fᬌn������XX34b"�1<��F���Q���`���>�4�]15j0p*��k�H���5l֛�(�����GN��0k'�p����f؄	�K�
�M��lV��r|aT{Ð8��a�2N:2jԄW�B#�&�E����/�݀���U|et�#�ge��\��J�0�3�$,�oڥ�LF0a�U|aT{Ð8��a�2K'?�5sgq�Y���!�fSk��ے��.gaBsdYQJҴa,�\"g=��)���q��m��6����,?b6q��i #eh;0+K�9���EG�9@��x��w�R���Y������y�W�̻��9��o�{�[.K���#g�_Ef����F̦vɔXs�n���A�a�M�ԭ?�;��4�u��^�.75��.�k�f��s����2�=4f��YG7b���00\��K�p�"�)\��m��6����,4ɴj�_�5��������St\(ؠ!#F�]�2p��f�,���f]�e��M��&��(:�Q�z��2dVm�Q�����pA�d�,���Q���^�r6c&�<.b�,ݥ��h�m�QѬ
2���͊^�Z�������ۂ��M�|� f�yϔ���,g;4��C#&Y�N�e�d���}9�a��\g-6��1��S�]!��rR��l�cb�ƫq+6}d�13�[K�*�yn8��sf=7��]�̵t�&�+��ȰQ�,�si��
4��g�B���o����A�����r�k3�{�f��j.Q5I{�v���\�]��n�|�58'��d���_�S}p^�lĤ҉���xKf!�s!.�.?E�,c2��ŧf�b<]@��&"S�fsKi�	�\��bKP��n��������u��j4f�,G71�ѐ�A����eFMV펹Y�w^�`��[@��%`2w���fb<�nl̴�+����Hx���$�޶�9p����܅�|WFM����Y��Ҕ����sBPj
9q�q����u��Q���|�X:lnmz^���s��O��'ݩ��9�M���z2)r����H�I6�c��r5p̬�3pR[Ϣ��\3T{�fm��2L!N3gO4�Յ�p���k�\H��Y4W*	jkw�]k3S�&C1dR��j܍)P�X�
��ͤR��ā�a��2_�f	�ͽ����փ21�v7���I�r5`j4�5aj��{}N-9d�T��p~�����I�}m͜+tcrj�
sY3����81�-��u!S�o��y#&F�;��.�O��Uӑ�{�Ã��/�A����W_�Ԝ;G͛��VQ�0#V��ͦ׎3������R�^Éq~ف9<�7��_P/@7d�g�21�Kxq���Z���\	1��ͮF\t9p��
^��H~GZn�ֻ�A��D��z,� ��рA�֋P�a�r&s�S�Ŝ�w:��7��spA���g{1�ȋt���Hz�]��ڒ��ٺzl�.�����\52b����=�ؤ�����SAɁ���z7f̰9T$�f��b��W ��?N=���êq��$�A�گ#������Af�n4O���_��N���:ŸID��qg�:��]��5	u9�����ͳ9�M��'�4JRnn��{l-^0��ׯ�������8��ü8��a�
&!�Þ�q\绚6�d��w$A�EH&�s2�/G�:��}2�$E7/&&��s#�L��ϻ���j�l.̸�͹a�����	�s4���SMx�V�yP�o�h�Ʈ��,����AM���up I��j@	"eh��a�4�j���5���[��qCl����q*h!�ΧX�g�E�����������ѩY�s�
c���~��3�<��F��������r�ˎ&��5���A6a/�!��/��K|���fi-8a/
��(03Q&GLN͑�f`QN�����ۋ�rИAS5�����������e���Y�p�C��F��d�"?�>|�C��"�&-_ΛJ@��^hn��)>���`��!�q3����"�&��U��+��hҸ`��q�&�浽�ksh6S�����I�ݘ!�&	�/�40��e�B�w������k�(�,����4l�<O��!�L���i�,�勦��kN.ߴ8fb<^,�i��t9��d�/�\�������/�¥���s�J�x#�{b����+���1��ތ2��D9��l١i5Wi!]�b�dC��B�G&Y�@��3�i��f�6�̪�D������O��V3�l���F�&5�j��i=�{)�Aӆ��ʣY}5Y9���d�C��kCݜ���m%��i���
�^x���u��&��
fnh"�V����
�����I��T�M�Η�,dYN�_�k����Z,�$k^�f��\O��m�=�%f�IM\���<�? ��"��M*�f���0����7dދa�B�j�w��h_�S~ج��T%1�【�d�p�Ok{�9��d�n��A��o+��=f���lVL�(2d��91x��v���e��a-3��*o�MI�������A3в\ҷ;�h��0f:�bcsW"{z%�\P1pu Xlh�d�&�����ĘQy����v�-�5]�C����� �e��٭�Z>�-G2)P'��y�� ΓL9��M�.�+'FP����E���>���d��[�c�,4���*��V�9��.Ws�'K�,���38i�Ɨ˹��L�=ľ���mBŵ�f�t���F^"1�96��FL��n���.�-�t�^KDM��f�fb���._�`t2�7z�q����.0�d1��C�J�d�1���^��Jŋ��S�+��B��{ �h�?��1�&R���L)�ĀI))������r9�4�]�x���;L$˛��Mr2�Z�����=Y��،:dڴ5^k�d��+|�S~��6s
�Q����W�b���
���j���[HFL��rV8���;�f s�/L3l6���r�!ڽ1��`*�Ĉ�C�@�&��9��r6���m�M�%�Il�a+`K@�ڭ�����m����,,�VZ~s�$��������Y^ϝ ����k�F��6l*l�s���P�,ݬL���͂r!�)��f�9�f�X��në[��S0�,�]8�D��!��kXʗ�y�S��
L��!sR��S$Z?5�vB"9d���]����k�y��pȤq� 0I���n�W�3���-��_��%�h�<6f�ȩ�="�+�sm��71v����r7��Q��su2W]�a�1叱t�td5�^�7=��SVN�k�f9�Ǧ���s��34�/5	��͂���
pn�2LA�&	*/?�,��r�W��!g��hV�M|�{�6�s�P�"s�d�"�Y�T��4^�;�&5�6q�Ku��yӽ��Ρm��ȩ�p��Q}�Ɍ�p�L���0p���#��m	�-�b����^���_�4S|������7Í1��
v��V9	 �Q`b��}g�_;47����U�-\���s��Y ��r5g�ڸIB��D�
�w���]��K�ЙVo�M\�4��禥9T�-1���������b]��)�������7��4k{�.6p���cL�&��FL�*�9i���,4h2�3kc&�k����f���Q�u�L
��\��:-W�E΢<.op����d嫾��+�9o�T�!3�J0��6��fm�˶��L�}6b:D���<0��f�T����bFL���$���4^�
�'�)5Y����6)-?0��4�qC 6þ46�JN\9��UuS��5'{<ʰa�T�\k���//4�k�X�d*ݒQ��ȷMG]�U����ƍ�s'=�?5W��e���wB^�D=91�[{2jN��+�k�vBCWן��LL�f�P���\	6r���5�,s3b̴�S��m�e��I`z���9P��æ=Gs�m����П�z3�L6f� �~��9��<�Jԣ᲌6)��K�z��7w�L�֡<a����9!���k���͕R����}m���.�b�鲘֞L��C�r��|��vUA��g��&���ʒI���Ws��i����4��{m���$���bԜ�n��z2j����\��QL���x7Y�W�%O���w���w#���tjt�9�՜��~��W�Z�GC��[9Rϗ��M�F�sA�9e��f~'����l?1����9e�M��|-�İx��,���ɨY��rR�M�}�݌��o_3`�ob.�8���EL�M��g(3	�E��+c���:��TA_�ͬ]J7O&���p�,5-�e��'%^��.'���O9/ Sc�34d����� _�����݈�Z�p�9��$`o���q�j��)��M�w�`�$�՘!3`���cf�c{���0M��w�Iv�Ŭߠ�H�f�/�K8�R6����_�g���U���'nds?����fQ��SY��l`	u7������f���WC�����p$�I�QI�������k�F������e�e�~?3d���� rĤ�3<!c&!ȵ_���L�2c��MDV7�^1/w3RV���)�&!���d\{����j��*���v�%b/51	���
̡�M���z�I��fc�㵛G_4b<K��+�w ��W��W�3$N�%�$ڲa3�%����ڷy0	&� 9��&A��/�E|���>NȐIPl�q�X/��N7�M۾�fa;Z���IM���΋�ө's�Ō-	�������Φ%?$,l+XMB�5^���ٽ���MSty��W$���4'g��hnK�6s�n~Ib.r�$��C�6'N�|܀����3��?ꉋ�a�� �(߸1q�sܝ�m���.?8��k&P��%�	5gq�A�I�W�L�ڋh��<��9�99	��x���}.Dl>M9����"���Mkq뵎dj��O�Mp�x�|��i8E�rN�Oxn�M���"���j�2 sxMx>�Ʃ����|O��b��Q���VSLQW����1SX�掯�J%��ib�G󚥿�F�m=���"t	��#GM��`֑��� �\�������➱����f�I�M����Q}�7lr���`�fn��:����d��Kr���	�������ǂK�q�J�[��$8~&c�C�Yr���Wf���	�WG�4qj�'8�V[��<�^�$���1����5���5ZAk�N*�s�<���4�@��_ț'C&Q~���8"���%�a��5f�,�M����U_J��9	��+1	n�D��vZ7l1���'�)�[o-f�'�7dV�2��u���A��O���G�o�0b�/���}ƶL���݈��z�A�9J�V�����6`�/�0�Y��73E��/��Q���)�<��8�&�E�t��fF�3���O8j.�5×�u2���n�ڌ�űؚ������^�SKL-7��ե|�`�l
M��]`��.?�w7+'�/+0l�$����Y�w�Ax� �8i��GL���dΕ�����وA���f��)'s4��
���͙���7'p��Ű��YцR8+���I�����[��L����b�k�|�J3	�{�B�W ��|�C3���.�era%����qc�c�5���7D&	H�6s@c����4j2�<�fbt����4�ͅ�2�|Q�Q�P���6b�䈙��S<���c����v!Z�`Ĵ�+�~��d[>kg�
s��˷�;�mn�R���������,����6��]�p�Tf8�/�l�\s1m�ag=�;����.��G4nԜ��"Q��S��hbl]bW��j6w�d�=��L���G�2-7:�n1Ԭ@7�o�U?��*�@[�4�Y`�}qE˼�P����b��x���S"��M��i����fl���w�*7l�:��i����c�O���ES����A�6��7#'��ׯ�1k�Ro��ְ���$�_���yȨ�/D�5�~������c�z/� �vd�$�o�dH{�c�9ѫ�d��2��Ф��G%��;~۫�d���d��S_�FΒ�#��/h�EKnf�72R���L.?>4	�7�� W~�oLU����fӉ�3�L�S�h��L5�<}V7h���,@��7uj�mќ�bZm6\n"َ�i��Ws�6+&�j1��L��G�jVz�"3�m5\��T��E�֯��5)�/��������Y[6h
�ݘq�|���6��T���$)|���18^I3����/�# �`0�G&�~s�vd���Q� 	�݈6�j��Jދj�4��D&Qf�����Ǵ�j�3�8I�%�FM�/�rV�&{/g=��+&�x��p��=2�B0i	(A�m�:��>\ֱ!tj��YS3c13��e��0�Λ(D�_d�ۿ���6�����/�55�ګ�&Χ���X�l���b��,��tZ(��	���ჃAlڠ�u|�YxĨi�И9��{��MT=�y���X~,�[�fcp�w���5���c3����Ͳ]o2rB�*vZ�o�(��!4<��U�Es37���.��*�(L5�r]nl�e�j.�!�f��7�n�T��5��[ф�<ɢ����f��Y
p¤��6�����L�����[U��f�ڕ$�$Մ�*,�܏��^�	ւ{�T����f��Y�����ͭ�e)&����Ŷ�W�ґ�jY�.8f�@U8dR��mrٚ�a�
�����a#���W�CKS�H�:�6�&�6< �F����YM5k��t���Օ_�Ǚ��C�f�,s3p�,��a0�ELsE�7Kt�n��=n"'M6��	3fm�d���|���pج�2K��Ye.b�,9�dج����(����R�pA�f����0�u"��۠����g6#.9�'3�{�v;3�=z.kv���t}/�pAw��+-������|D/�$�m���9�_,9`ؘ�Z��
\�{�Մ���	߶a�e�/ȫ��-��-to�� �1�U��PcFt?�"01k�e�0nm��`��>.�E�@��z���8wr�v#�6D�}]@r.��5ݣ�@tD�#z���[�"�ha]��\�5�L�q��YѠ)
nEfyndq.�urZ|tS"/9���Ldn�BxE�D�*<��@D_���ip�E̚�Q��':.����M�`	�M19B��LT��#��.D8�GX������/.b�d�)!F�*��2l�Հs堉�UxՁ�� o��=��_ltĆ
�ˉKh"Í��!r�Ɇ�آ]�6����^mc�r޵��F�P6\�%������nU2�=�wV�#R���
�Gނ�$LuԄI���7����L%���20���\'&"�,�[����,��21g22������:�̜=��&��W�=Z@����Y��Lb�Ī��*�Y)3c5�Z��AJ�D'#16Bɹ�\Ȑ���,�#ˍ�\h&	�!�Β~���ѨI�ѫpBU��qy���f����z!A3�����	%>�1Su�	Yr��td2wzcf�$�X�{)��@M��0�!J��6G�<*���
�/O�dݼ����RZ
p��fݷ���1p���|�ݵ3��6+\��ĸ�sO7�NCD2ۀa�f�nj��.p�(�����И	���f	݅��NL.��3��8��$�N�5VC�͢��:6�}Bs|�p�B2���| s�HYDã����̺/��s�ã^l��p�E�0J��5�xG�0�����%��`p��!�"N�b	g�L�n9��(��]vrԼ�Rm��;U٨���E*D���f�;	f��nL�·:����T,u!s��Q#�'$x���ވ���&jYIN�ͦ�Ǧ��ASЧf�����f��I�����)h\�[�q9��d!�UZVd%ַ�^��T�l�gL�
&����,j�A���o�5I0Y�%��k�X�0���u�T��IĈV�2[�Y�����`��7�y������M_1h*��,�#و,&�G�]�'��=ja��Bv�ͬ�>1a����<n��#��ѧ��me�d�s�4r�b%���Q��!�$aA�)�ܖ�ʃ)p/���V/ɻH�`s8MV����l�2]���@}��;�(ظ��R�:E(�~]�l�İa�?9��-�.18�P1�1�8�o �Ag�"����˩K�͒��&\����1sT/ɢ�Q�9ݬC�of���s+K�U�s�՘9܄�N��&�,���U�:4��Q�21nf��6���݅b������i�e��t��U#f?�>��e��0ň��>7�osgj�H'D��%�_�0��h�4uח�幚W�d����T�Y�`�e:����]��^�\�}��_�^���@6�t���s��Y}2��Huj�\��.Z4�S怴�k�f�V�h�#g�gB�l!\�d�,�e}�D++~��#�;��SaI�fX&��Wn�벃���|)�^��#�6�X��
=�R3s�$��w�����?]��,hr��$^�e�fY�Y���Ϥ�y �FM²����qm�
���s������F���}5r~�\ln���,�������嘙�ŶN+�b�nJL��ĸyX1k'b]�O�*n^�(h��;��Y�+m��������ʆM�s�yU���X���p��[�$���2Ynˣ-[z���}���F@���V�29���e�c0C��QA�B������=5<��$���݃�15�D�rY�eƦ�;	^r��,4qB33 r�U�E���-��_nb��ʱ��Ѭ+�M���r��+t����n��Uæ�m�]3�鎯����-T�*,s3+DL����Ԡ{Q�!�7�s@]�k�9�Mįɭ�SoVZ����.�wٗ�uɻ	S�(��|��w�8W�	��@y�$����0/<���☿Xݳ V�|Y	5h��d��B���t#f�t�g��'��N��z�a�.�s"��n]ϐ�pmɈ��s�Y�b.{���s&-���L3h�Y��Kjti����^S�Y��t�}�$�23���}I��Z9d��s�'��"ll���p9�n�3��d��Zh>n�\���pi@s����jR��d���d�ٺ����uͫ��5Rs�ֵ�'格�b�$��,_8�K���0��<�JI9��:ܒE����V�<3�G&i�O�YyPES���F؈A�f���M��Ǒ�⺜��<�75���?O�תI �@�J&Y���,�e(�@�6s�.0Ip f���,+��Jmtΰ$)nٲ�������lnw�w�z�o#<{�e/�9(V�L��N�C!2� 2��+p-ܠ6�Ir�"3�sΛ)���L8�#��J��	*�>Vןs3�jm��  �=��J�m!����t3�%'�neG�%�������z���+�꛸�����輏hV�2=~eˁ�{؏���V���M������hW�ŗ�3����Šf�������������xb�Kf(�j6�{�\�/:#�v o�p�\�P�[Q7'٭<ĊYVSJ*H�<a�du��m'�0O�z1rFq9�����/��:�1SmS����!��Y�k�ex�k��I��j�Y�u=��m-ds�> �ـ�d�@������u+������4��k~(#�X����Ή����⹉�b5'�4����&b]��-�s̐3<����.n�[2n�k��3ov{6�*ds�?��i��3Z�؂f
�I�r7�<����������.��.2I25���Z�h�k��d���z��͐�hKfjJ�6d�_h�\��W���1�n|sP���kͼiz�G��u5���LBڲ]W0# 6��2諸9�ь1�E*\�Ml�V�&�g���u��mDB���]x��"9,�Q�,DsCج�-C���|�Z�ͫ�#&�(�̕�s���&j!���me���?��cY�+��k�s�wg��$3�\���2s0��bذ9��Yh��d��	�^�`
e���,�����t&P�d�7�X����̩����"�e����%���ov]N�zu�<8����Y�W3+���D-̾>вG���M�b��Ӳs_ɜan��/*5ID+<��lne7�&	��
�p�\�l�htn�q���r���'	7pbtRs|_��]���uY�C��[�u[!n�����Xrq ̝_ԋfɐI�W���V<�6W��/501uw��������a����c��LV�[1�s���s�d��1c檻���iz5n��,�$1�������t�$�#��hέG����]'9�0k*��n�IB����	���ȅ��Wb�q!�	[7/;<�yoX0k8^�6�Z��"Pہ�
�/O�dYz��ڂ�+�`�q�Ƈ���􈁳�/�������Ћ�t8|���W�Y`�\ϥ��Π���
��ůf�����^���*���2��Jn��duח��� q�D�+>^���5rΠ����i��-Dw��Cd��98���0d��!j�ߠb噻��6�>��u�2StYÁ�m�.��:l`X|�cSb�Y^�fE�Q�Z2K�Hi�n�L��su�,�?��Q�lF���ma�A�p��#�I:���\�u�2]hf����y��f����4������Y�sb�A���
܃��:c��)uYw6l�lY�K�=�hX�u��l���S���.w5_r���p.�8J�0���2G���Z5�������vnt�i�R�".f5���'T�«��}#��z��s5b6�����͂w�]	8Q3<.7n�Z3��c�/h��SSN�q������#������B3h�l{��څ�P�S��f�o���
7���YN��FﾛM��Sr@�l##ݹ}]6l�D-̪�Y���<Ƞ��ĈĖs��ʙr6E:E���� T�~y�$k�h�4����~!\��]"l�Ԟ{p��w@�<4��q�\7j��3�����?W���:4n.�a��X��s]��uC��u$��p��U����(N��l�2�ft]܄B��^���^�f�~-��ݽE#G8!R��(��@��-ԜeW���C�ub�Qݺ(�Ь���Y���fܰA͡
�8h��/"wK������Ph�l��[�t�5��뺙�Vjۺ�Y��p㫢���nٟ����ac�m� O�aCˤ@�ԭ�	|#�}�-�n��s�%ʦcy�ݨY��{.6�|��#�&Y�<�qy�+��e3u��p��9��忊��Zi4�n���&O���n�����3QN���ZV�1UKJ�5n��
��ʓMM�˫*�-�;�0��u[�5"�F���7�4Zׯ�V�f��6W')�>�<򩹒��df�8ɺ뼩�pC��&_�+���X�^ε6m�,���
�
p.�ɺs㬹�x5�hZ33`�L��k�~�O����"��`��A2n*_��ʞt�*�L��ͱsCī���hy��X���[T`��]o�7�f����6#�巑ky.�Be)���!\͉���`c56vW�y�?��L-����4h��r_d�tu�������[�{�뤦���gѿ:�n���{�[���=Y�uu�r0��U\��N5�l�}+��&�-�f�T8\���;������$�J�_b����^l�0?tZ�a�rpSY�������ɺ����F����́c#gƁ<I���@�rX�P�;�?��e"fYM(A� ��I���{��vB/�'%3D�g+9�g�Vn����'�T���^��uh�cy�9��Y��Y:{��w��Y�.&D��^��uCGL�.�j��b�HnJK�y$���-ve����9��K�L�/1��߆�&���nt�B�nݶD�A�Ԋ�����E�csҜV�Y�9�:3'��^-8<4��+�TAЈ	1�*l17UN�CF�2h�Zf�$�ν�F��O�b�J��!C���ԭ�!��A�M%Ċ/G9rĘ9 �I�q�����	�&���������u�ꐴ�㺜�uſ�V35n�Õ~ٮ�Z�j�"4�6�AL lB̵Z���j���w�@3�'ӟ�dVruW�ME�ڳ9��tc1���v�l:�=6�4���ß�;�S׭<7`�,/7�*i�����}\0l"�e����ZO1狘����k���@S��F͂��̿pĄ�n}���;e�K��n�e}����\�{`ƙ�3�VZF�G�x6�����s⛩���]M�����1E�R�osz�C�[��r��YڇK7Kqa�,_����s�Z��C�*�9}԰i��Κ-�m�H��ԭ�"4g����hu�Wb�j̨A�ȓƟ�r���#�����W��'U[�[���w�&ZY���usm�@r��p���	�x��.��r�t5pbI���j�/0���_��.%1KKLZȜ�W�ͱVI��9��8_�����v1���N��)gC]%��}\�dȘ��sTa�I6#�K�.���pn�ʘ!S�#zz8+����q�׺��&���N���V�M[�W_�ˎ5�o�!�&�,2n6�x�Բ�^�[_-910����<b]Ω�L3�p����3u�l�\9�@�)��v�����&Y�F3���� r��98�I�Y\`��r>��쮝�
��c��͑��a�^��>�q�������WC���B�枯8Ip����;txߨ�D�Z��斻	��e��C;�Kg&駘���.
9j��	���zD�/��Y1��ãfl��p�E�.J�����v�b�$�?��'�E�&z�(Sz�I5�`��9��KϪ́{�ɰI�t���lf��u�A��o&��-x��1�,F7�n9.�bVl����dz7�w3�nڠu;T��
܄����6��j��
a�~��K#gsrh^����5�������	�<E�a7d�"[L)4s2���?���a�/Ës4-;4a���G����4p�#�S���!(1a�{\7G6�%�
3Z����5n83��+p��9l�)�ق̝](7�&ƺ�3�������y>5���a�nF]8��0�r�;I6.��ڋ�c��S7�}6f�Yk�t����!��0խP7p-#Eҷej�:U���ϝ�����L_�JL�ч��I�]��۪/4�D�Q��1u��&Вy��[�9�C8Ic��\�L���=8��lpm�D�ˈ[��0��O��� ���?%�ߕ�4+��~��t��J-�Vw������n�`�n�-�7-50rR������R��M��YX�����Tœ�@5��i�e�[`͜GgZR�(uc�l�X�����l���Z.p�TD�Y�5X�u��$�Us9ԐY���!�.���J���	Wz8pn�smܸAS\_��ւ��Ȑ	S݂}��Z��L�E(�4��pQ-0b�$#,��C:5��'�}�虶1:�lf���&�&b]�a),��_�rA�FN��G������tu�İ΅f�oT�����P�4N�`�Rx����a=�$�'�e�)9���O��t�ܬ;01�-�M����R&,D��d\�f܄'��:0�f�T�[ll�,^8~nR�Vx�!����I&D�[*rV��]�p���>mgu`M���2[&I��1�ΙCNĺN��|2�	S�(T�D�,��|�D*��v�����&Y@VH=�pY1�8Wyy.)8���Y�B2�+`�\% f&�
?,�y������g�2X�����asgo��/<�v�\�M\!������c����٠����>["�p����ͦ��k��\��,�+�����_�;�o\L�b|_���͒)���
>� 8�k�N7�|+5E'9���v�^N
&/d���`����٣f�l��Τ�k�^˗���+uG�z.��r��&��r8��T��9�K7k�Lb$�4�}W�M��̻M�9Բ�Hz�b�M��{�b���!s	,�ú�p����IA�M��H�b��)�4����b6�Q�uW{Y�Y�j���>k~2��j-w3]xTmu�51���z.K4�\���)Ow5�R�E8b��.�b�3p.Қ�1��&i�M=��Eͺ����驲T64���;�4K�Mҙ��԰��عd�$�h̠Qs��d�qs6���"���S�M�ઉX�)�j��ǅ_�!r�3x)���9��`<��X���R���m���ܚ�YH�uKPÆ��.f��LJ�Ksҳ9��8_�{(�s@\j1 Hf��|ae3rԺ5�꾒ِ�$���q�͆|6Q����z��h�G1�<�<�y��� ���i�f��N�/�E�xd[0���I��Q�f�Z'4r&�r|�Jȉ��M.����]�U�Z��DF���1��S��r�����L-T�	��@	B�'L���i�� ����6��$O��,��,���b��3��Z�ЗnQ��;l܈���s�?��l�L�&8o��0Ќ3pB�n�l��E�*4���.�ཁet��	W�����j�ף��rr�l���l��/^��T[�L�WtŲ^H�ͅ����Zl���s�\�#?Y��>��Y���H��ףgEVlY/B7���Hssp��r2�Ȝ.�����Z��U2�d��C&��pw٪�s�1d1�kM�}Ֆ+�S�����nbY~f�,�˰nnj�)���d�����ly�9ਹ�f�D-L��e������*�Y8�,6�T-�4а�T�[%ݜ&�鬰�Lhν�f)�:�P΀�p�K��~>�/]�ץp��LGv����'�8��Fsp� �8�i��L�ml��YC7`k%��puq�0Q�������S
W������lL���f��>f�D��~>�°��W`Є)�f��c���b�N�ꄩp!��`V𵋁�HuK�
n
�F�$�zG�� ��K����G�51����1�A7j����Y'5n�y9l�6�	W�o���eV���/%0�K9`b�����vA�%�b2��ۥF�6����I��z���1s�-�)h~��sX�i�c�ШyP6-�*��v�����&Y@��������b���B�S{�,~3dp�,�W����l_���[Nd��Y&nNK6�j&][��%g��:��%��6���3����u:L��[-\��b�r�$cB���Z��k{��-�G���3��S��pڝ=KM�3�s/�%æn�P1k�FL"��lz�\�ˍ�R(�̇�zpF�4���{�֍�ʻ1���'c��i���++ga]��t��Xy�Y�{K��0�YZ��gSI!G��p%�-p)p�pi!kى3����Q���g5��N���=�͘l'b�Yvr6-g���	Q޵l��U1C�.�[;��&Ι��&�<4���3~�s0W�BL�:7+�8=~$��R�*�-�m6C)1W�-��AӅp�`3�$#F��=N��}R���s_%s�c
G�{X�\-���&I��?�݀��QS��W_ `"fxY'1鍟_����3d�1�2��/��~����vS'��7�&iq��{�fs����(�g��&g)-"91�.�*6���M!��%��{Y��Ĥ��+}WKN�kM�,37f�����
75��sV�@ݚ.���yk�72gɦ�;�$q�\�ã�3���@�RX��1a�q��ܦ�['8p�3h���vdȄ����:nhm�$}�T��u+��/�11�1r� S�~��۷�b�$�9�u[��.ra����>�Yp̄+F$�-�(�̉��O0�������+���Y�j7�E�H�
��0NS���<웩~���k��M-n��RZl`И�Z�2q���fwI��d6�n�8�-xG��2���P��Y��f -�k���	���&.~6r��iD�8�L̠y��:��
l�bЀ)L�P�`��u9��̈́+F���nί�m���"N�@mJ*H�<a���.�����[�a��=���KfwA\�Vi-j�Q����D`SDs@?\_1f�d��pY:b�3e�&d
���q�4W����In���2���".�E�f��~)<����.�����-	3��N�5[���(���/\VhH6�i5�Q� s(]&��MJ�W�������Ѳ.{xS���G�SY��k5�l܄���]���0�r����1s_����'�ʍ�©���g#fH��J�R�Rl����uj��I��B#����s����Z�2�]W/���8>�,$��!j̸��[31fЬ#1/W�,\_0����
p���q�M��jvj�1�p�\��{�gO.�幎+����)���x�pbH).p7�V2U��.5�s����!nu�ى2���k���0O�Ph��7~��_Z�� Sxo7~b�1Q��g�z��S�&L1.��YV��0Pь.�wB3�*<�o��_N<E�{�&�,0bиI���,�%����Y��]���>6>x��0�t�S��Ҟ�d�c8{0!�B�T�A#Fι�����e���{<�������9���l�1V��X^Z��u���-��&���Ud3�2E/4������BE���� T�~y�$��R0��0��8Y�~+9��&,��Gw>35�a���\vg��	����K}�ݗ>ᚙ5]��n!WN-tsV��UQ����h��2qs2�!Ӆ+�������$���'��-g���e�^+�f��m���ͳY�u��N����*/�%��,�%�&L1�K�-X���$[o�K�Jc�z���d�^�գ��`R�z�º��N�ʪ�8�c��qsB%c,��}sej��XC4#l5j�1�pY/���ޅ�h��	p�Q��ɦf//9��M����#�ͅ~±!���g��%U�[�k)�<����������^�
Ũ9D,�E}b|]��8�n�B0p�\B7A��I��f�+�f�%�Z|K�r6��1�s�?��84f"�eީ�-�us�K����6�2�Yߨ�xI6tX sg��!SXjk����:�	S�q�i9fԨ1�<�$�Tx��,�u[fj��I��4yf8Q���˲8�yƵ��J4o�{�bԺL�el-��vS8=¹s�����hb�9���m�5��5T��>V��u�������!LD�Tx��Y��,�OL ����)6)���wf%�l:)ٺ=���_n����Y�Y���8�M�bld�>�řɡ�b�Cu�B9$1鈈�e��3�X�����巩����b-�X���T���'�ڊ�0`Y�ռ�0ňƖ5>-�M.�Z��"Pہ�
�/O�dY��N?�ps��p�\�ku�S{Vr���p�K�̄��e��a�h���X�%�Ư3����C��Bf]�QN泜��7&�L���(f@�L-�Ԗ��e!'ə%�f&s8$�"�G0j�����A����=�ψu�ߺ/��gt�P���͐a��S�;[N�{x����� e�ߦFN��h�	�)�&�厈�#gS�殐I	��g��d�_�%	���,�+謑������i�f�����M)\���#'����J�6nr��]�����֌2�ky�Dqd���;t&�I��
'I~E��ccY��gQ�TQ�n�z,�uS�&�_�������ͩ���t\��=Q�����<�&�����h̬=0�7'�*�Y+��������`�B�B0���C?�39raF���Hksjݑ�F�`\���I�rМ��pd���Zn+f�ᤖ���]��9��
%f��U$s�m�&Ƒ�kf=��v9q֮���_W5r��)B_����ySR�� ��"ް��̂�Ƈ�G����Bp�/�-�h�D-̾�eb6}+ܐ��p����.�*�f���Z(�Ux��l�[%A/Z�&��}��`�������^�`�TxZBlN��ǋ��^�U�:E����l�/(8aJ
�as������
��w!���mYb�䴩鏦|E��S�f؏fy��5�:�qs?6�1�[f�������9�XtߏW8a�q�ĬO�g��[���>�7�(�
W��3c桶I��p@�6b�l�q2d��v��Wg��n�8R(ޝ`��쇕��� =�	�f�\�c���'�7��a�G0'R-T�	��@	B�'L����z���_�Su�����������3Z��p�_!Ǔ�f9�u��Ѿ@-��L9����wnԀ�S��&sګI���Y�W��!S�܍�"gu�Q|�`k����N�Y������)�_(溲��:�Q������)9KVM�%1ȸ!�۸�Z8�י�������^�t���2}q��\��	0n�1�=��3o�Q3�	�m�s�c���l7{�S3��4hF�j�$c����4���n�<�b��hМ_��*�q�0�r�G�m\6d��U_�s0dS�1�\Bs�g#&�n��mݜaW�vr�zE+����M���c��FʹvᓺY��4���^l�Yy6�-9dj��7"gn��k1�AsԬ�4f"�eީ��a�.�Mx����P�7��n���iS/逘͸Y�w�2�8��n��ud�«���S��-9	G"��� �Y�e��$�O�g^��Zx�,�b�<�Z�A%���v0f�D�˔\�f��r9_�	S�s�p'�S����5��RHJ���xQ߰�+���R��r����H��9.�0%Z���j�R��l�@�M�³��qg�8I���Yݬ�r[�D-̪/�j6��(Y[4኱��ab���,N5Ci4f�P��`s
�D��2B�s�Xȷs#���Z;1nn}!�1�䫱�8��:�hk+FL��,��6\Ws%�	S�H�\#2��K���BE���� T�~y�$k�h�N?�ps��p�X11��*�����9�R��L}�]8���
d﫡���I퇳��>M3AL���Moxi$����[��;�j!�Q ��K��h�ia��హs��2-|k~xI@�W��w�rf�,hU������&�D]���i����}/!6�g���:�1æ�eK9�4bRlN��?
��ALƅ����f���I�k�,���B�
7�恗�N��:�3�z����Y79�]��)xX8h��Xn��ˍ�N̺�/o����I	_��$Za<�>!�3f����9���kn�����|�:6dVb����M6l��
�s���S�r[����+Qv.��3�7Ѫ�OhVa#G�!rͦո�s����z^�A�
���[�r�e�f˅��Y39�>�O�1��9���ʭ����;�ؐӒƮ�a��G���7�F�Q��̊�{�zL�3��s��l�'Cjĺe�A6y�Ô~AX̏��g���ܬ�R;�i[�7w�� $S>Ŭ1l�D�+��YY97Q�3p0�ͅ��b�ȁ�b��Z�·�u��ɺ��(]������ϙ���AQN��g�	�	д�[-��o�a1��楽�oښ��p^,�s9�/nAЕ=mע%�:D�[�C�x'���,���;�-����B'��K�[�*�u�?1��\i3���ӿ�6���Gv����.�k��;��lbe�:��bW#綱����c��sH #N�"ԝe+q΍X�����E�xw�nM�8f�쓉��5X���U�"�e��ItR/ⷅ'}�}]���3���"N�@mJ*H�<a��i4@�*������^��
g+9�G�F�z�y���L,f��n!�Ͱ�\&������M�.�b��ኌ��;rϽ�uC�Q�[��/q9�밝(;�K3�UUe�j��L��~��r��9�{ɸ	���FG�/��,��y�\�8��Vl��p�E�.Z5[ofd�>��EC�,�C|��Qb�L��,o9d6-�-�u[�h.��s��$Y�p	��*�'��L���훴>7l�sY�gLP-ͥ�����nĺ��yt-1W�Lxң1�d�+��d�[�3�s���(\7K��I@fcdj�uX�{mf!W�,� W�����L�� &�4�sR�uX�nV��b9���e��٨Q�F6j�`�,�:����ޡUt�8��IƈRx��Y�-���d�A9b~�>fbT_�+����j�Z/nN�uޤ���Y�Ԭ�ZZX|U��jN41�3�0�`��48nV�Luf#��f��$[�j������:0O�(62�4	l���ά_�v�6uռMN~#�Z�s��	0���>���r@��M΢Y��]NK���p����H߃�5K ��@���9.ь=d�,�8��[n'S~����B�\�Z�=�&��&6���������{&F�v�!0l2m�z7+h��9݄�PLq4f�,�$/#n�ƌ����pB#�<E�Df�VM-3��s-oy�����FNQ=BaV��-�̡?\1��e�Y�n�gz�N'D��%�_�0������㝨W`�eN����"�������f&4.r�9h��Ĕ���we�$Y}�l���g���h/��M��+��ᔩ���TfV�RO"���\���#S�_`�k#Kb�o�;��FN��짛�:��4�p�X��] ϋu,�Γ�9.C�v�lx�B/5��3G��$J�\���)jo�@���������`���z�uX21:F�E�`qi�u��qc�	���}v�a�����AG���FLXb����
��"�vWG�)b�T������)B�.�����c1���7u����l��<�5���ދp�n MU}ݗ��#N��?uf�u�.8nV�L����7'�M�d�9�[�8���pw8Q��j�l�p����!xi�ص�` "nb�����I�p&R���ͬ۶h�$c����g�%!.˚ͥ�sD.1�Bs�胒Q�.Sv<̲rCFN�!���ąp��_Rpjݹb��N����H�ʪS�?��=�׺�l���x�,ll2QNw7'�C���x���rsјq'�ߎ��l��)u��8�^R�U�f�=��6Q��dǍ��x��	S0rn�nwt�B6[����q(�Rx��f��1��P��%����IZ��j�K�Lz38�1uC���X���Y6p6K��'��pň³�����<3�P'D��%�_�0�b�����S����`���S{VmE.�r=�굨��oc��-����ljI��qn<��H��K�)���,I����B��pGMD�g�j��VˊhVqѺ9a��:�'9��L��a=6Vүۢ��@my�'
����.36Ǯ�j!���kFF�6n�$��r?��AN�S�ʢ9D���z�@5�LW6Eխ�5'�I��v��n=����B^�;��1�.ƅh�9��-���f�_���L��n�0��"���a���r���l�t�t�D-,�.e7�b�9	���ѐgū3p��������d�B��M��ɩ�9��,�u�l������/���f���s!#�O�,�k�V�b8� ���B����X���e���&1���,3���炩���ŷxO�M����$s6�o@��쫘��]Z13�-�c���mBsgV�B#4h�Y7�L̜&f6��n2��G1��@¡+L�'��rQ`�$y����۹^j�ta!�<��*���,ݺ�q�O&F��9Գ�+�G(̪/��ą��ل+F�<��u�s��qBj;P�PA��	�, KHS}��s$]��x9��JN�s�#s]�<�����dԈqs�N߃d�u]���$��������TO�͈A���r�on��9]/x5��:nja_����Į�s�Pb�3j��G����d�G���
c�f�o�MҙH�[�Y��A��?ΙM��`sE+���_�;���J�Ef���8��U����b�b.�2]O3����?S�q��9ؘ1���� ��0s�j݁i!���-1a*��!��ٔr��#�[��,e3����N���P�&��amQ�I�X�E�2+F�B�u9Wv�Y�d��v��,/9�/&LDY�Wq�M�Y�lf���Sn7��F���YR��r�B9��a�ޤ����2���G��gԺe��/��&��W{���3�R#��v3SCF�11:-0n.���4��fAx�r��t��w����x�B�N������f�D��3�e�\@/zz2p��tI�S�qM����7���r\��^[�u3d=�,�����ά-o4��s��ul�YBK�e���o�.$7�Ǎ"��?g��#�uM/,2ǈ�G)��f4as����T3J�zm�������<�Yp��S�e��� ��pR�Oꍱ9��)��PX�c��Y�`Ԍ��q.���h&;s��{�d2�*4s�V�P�6h��F*�7��>1hb�Z���ِ1S�,��W�i����f����M������ʟ�h��)F$.9r��d�>��n.�5���R��b�qs$���f�3̄�����*3�����ͽ��ɪ��=>܂��0�L0�����6኱�Ьĉ�Lو)�le� ��̈́	S�q���K����Q
��Y/3{Ky����R&#��X���ip�W��8f��}!ja���f��'L1"�p̼̑����8!�(A� ��I֦� �.� �0 ���B�S{���t2-3'354�C���4n��h�q�٬��Y�АI��n�#s�Nb6p�46����vB�pѱY��by}I�ݢ#E�u7æ֭�񾒇z6Il��e�^/4pJ������d�&�iy�Yp�,���$���l�AR?#ՉqF�	�L��d���9̡9����jn���s��$Ssِ1�ۺ�� ���$faL"t�b�GMt�E��У��G�sS��7fo����$z6O�YhHn�
7�,=3��.���aƍ�Z�|����I8q0}й���C���V�Е�)\B���(0r�D-�~�Qs������j�E��S� mb�Gf������mɘY�W
M2����Z�)j�A�朂��vŨ}�-ߕ^�ӫ�`��y��#Kse6vR�>f
l<�B�f`0F������D-,~�'j�\��$GL�",9�l1�����'�%p���Ib/R���$�k��́3�g��ͺ��+�L����d�w�Z����p�9��I�s2��đSU�ug�B51��̂xP�s30�0e��X��"z2r�l�0s�dg�,�M_ݛ��v΅,�s@(j�a3�k$F�0�O6#7Ig"�t5'���&����_�جwU̫��pF���l�y��E�&b]�:1����d�Y���o�f��ऩukzT�9�c�r#���z��LZ91����$�j����-%ƥ9�l5q�P�>n�.����C$�S
��T+�s-��Zzb�<������s���Z��Es���&#&\��8ҷsS}\Zk��KK��S>Luj���cx�l1��41��TԸq�����L�=͏��B6�����W����t�13�aJ���C�9�ؘ���8!�(A� ��I3o�0����CfI-;8p��S{V���z�93����B��6pl���MF�(�D	��^��Hf���Wa+\�ŉ����Y�6��6A���x6��q��.��bn�A���3��"X��@��J���v�Xjp��W4�;��AN)<q��#lq�I�@�Fj��ʟ�dj�2==�29��Sw��c/	]��_��םL��q����g�B3�E1�o���Y�뽔ݠq���y����v0b�� �fg2�&|;�fy����1F�l�����j�)*��Fdv1)��۴�����/��
_2��:��b�Y��@�ASc\�嵎n�9b����K�и8�T��\�d�G#Sx��'��-�G�J��fWh�d�}����u)�O3��N�'�z^��]���Mq �Q�"�'Y��l�6�v�.G6�S���ĈV���l�17C��#�
��Ĉ�#��a� fS`���S8~^�1�rb�{c��s��nf�3�����@�yz𶯅���E�̀W��� �:���Zg"�Yԫ&����Z�S#�.�����\�����c`�\.K�M
qBj;P�PA��	�, +�\� �����X���x+9�簼$W�rЬń&��F�3@��!:���qsN���l�(0s�^Z����-l��	� ���+��l�ɀI򙌚c��I�f�8n�:�����B�fe��9S*���̬k1d�,l�e�nb�yX\h1.�!�P����)��R+s�Yp�X�Tx����$V�.�{��`��2Θ9�Ԉ�j��@u��ܰ�lj��!�͜�h�f�؜Y�C��p�8L�'7'-����ws�~#q��Q2l��J����~x>��<bR 9���GN�q\#7��u���q��磙���fY/�ê1I-93j�q��Z�Z�Q��u&Wf�7�F�J�)���Y�6O&F27K9n�p5l"�e6�9y�����`Κ���\�4G�0� 3rr�@�¿���QQ�<ܪ��(��7C��@���{O̦��fv4OI7n
j�0fAN>����<V�`]!�=D�'fЈI�<6xN�����ʢ�Ā[�p���i�FL-�sL�`������e�k�,\{6�PΝ&cf�-E8����EH_��	C�"N�@mJ*H�<a����fmO�v�����Ԟ�{��2\a�����3��Z(��C���沞.'�%��z��O���3�_�0dj��C2��&��U<��S6jZ�u`�fp���~�'��_Ý���u���`s��I�-��}5�\x"]x���Ņ&��9N�n�#j.��sb̸I���J]�u�X�X����<1�8g���d�p7k��[��A�&���\�G�&ja�s�����#&\1y'݁����5;�7q�f3(8�.$9Ee0l��Ձ3�%���kt=ݜ��b9[�Y2��:��b�Y7�ﲫ1�	3���Y"GL���Fo��S���f���!S�����s��_��b��f�W�d��e��''b]��S��ƶ�S�I��C�U^�`а)�3 p�X�dẳY�G�27S#,�G0�S���ĈV8����'�H��"��a� fS`���ET8.�a�����ƞ���V!|�ܗ��-��@�i�QzZ�s��9��6Fؗ�����e ZFK�ٓ����Z�SS�9�/2f��a�N�pCg��0*��v�����&Y@�1}��<Ĝ����g+9��l�)���3SC�r7��*�@�B�x��޲3(��鰀���%��ht��˛4��w{Wv(Q
�G3k��l��@�Y�!�r[b���/511��Y��<Pkfq�8�p	�9hʑ���$�99������PQ�f`h1b��w�ݪC�J�XZtd6z�X�`��	�+���=��	Gz2\V�&�Ag����
�t{bN�p^ȋi#��
9j���r�6���g&a�P���/W7ى����͞7r��.E2l�,�B���͓h��a���1a"�2=���dԬe�u[��~��&����v��뎦 ��jf�>f
�Q�cߎ3=�8j�&�sI,S0`b(y�Ŝ�Y2`*��Q��ɘ�nQ����<�c欭��&�<��&W����Z����>�rɨ��2��W��8qఉZ�1�J�j�� 2aJ��X�FL���AD�`a�L�&Kt�<
8nֱ�a47�����
/�c�Ư4n�D+\J��,�w$}���Y\�kMԀ��bζe�����if j�p
�ϻ�4s�<f��HuG�f1B>l/2G�Z�)�vT-��Yw8)Q�WE�91���ύ��ϧ��S/L1\�\E2ř˱��Z�	W�6s�k�&�k��e����87(F��92r
M���xd8���fn��V�&ja��������S�pň�C5��3�4�G��n.�=5dN�B�U�9�ĉV�����a&����l��UsSyvT-�Uvs3�h���9�6��N��������G���ٿ�b�d'N��6I�p>�F�5	_��Y���g� 읹�n��Zg�lqH6s՗��8&�y�j�����Z�2��uP�N�bD����ll��a�BE���� T�~y�$���`�F7�\8p��S{����.�e��B�<�R�2.��� 6g��{�Ñ��77����\h��Yt�M��u��X�ȑ�NO��{���,��L�M��5�ʊ_��EyR-9d؄%��È�n�`�e뷠-@�a�M�m3��}9�̸���as���aF�ԉ9n^7�Ͱl�>�ρ�bmbү���`6B����+�3O�(�Z�����t�Z��\Y�'쾚d�(��¿�Ŝ�r�a�N�Y��3�&�M��d�NK�jC����h���5�\ͩ���wN�
7���O�˺xظY�bF��3sj.m7^�$'��r^�b�dVH[�tה�8'>8I�O�5h��up�������I�	�rd���i�(�-u0j;'�7qp̬�Z��?��P�&�����k������_�8�������k6x�P�x��as��T6aJ/����Q�j�ɲ .7��k��-��p�u[8Vz��&<un��b�Ac�z%���.f�����I�_Bl(nNb0��
���VƩ�^h����u�?8l�e5.�)y�-�Cǚ�j��qBj;P�PA��	�, f��.`�иn�ȁsȒS{.L3d�!���h���sӗϺ�����-�bи9u���'��5^�r�V��U>�-��ninV�I��a ͚F/8l
co�Sqsge��m�b��a��T��9t�q8K/�\0l�����}k����Y/���J2����z�2��Hu�g�ѡFMҿ(u7��p�!��nܿ�.�격�j��,�n�����pԜѫef��O����B|�@m��0�X2lȬ����:2�]�ۺ��ʈ�4n�lLL�=���cr� �LY���ſ�l��������I:q�Y���׮:p@޼�GZ~	��
���NN���qgͬ#���Mob�X�ܽZw˶j[��H�f���T�Weέ�ͮ�7�FM�o�Y�ƶ�����fR���k�;T��Ʈ�*m�S�E�[Q9�X7C��zĺ��J��u>��I�������9��ܕ�K��R��;�6\/ bN�huЈI�����jʁ�`���`��a+��j�ຟa]�p.�C�
L��랜�h�FL-[v�u	,C8�oc�
\���ں�^��"Pہ�
�/O�dY����幮�?�A�"�g<=kf�Y52�f�ZL`1Ǖ��e�֯��s!-1]6p�K�10wM�"Z�r�U���m�/�&�Z�lm؈9���y�6l�l���e�,�s���p�$��j��j���n�*l���f��ۺ/�p.�����-�����nM"��f��r�W�L�uݻ���М|7wp��4b�%��O&I��>��;��T89��Y��5�@ˍ��z$N5ˊo+|}�H�Y3aJ~.�uesTWߞ��� ����_�A��SU[Zp�9k,')���Q�f�9N��a'��m��N���Vkn�D]�r�$鶪K���od�7�>�KV�Ѳ��KЍ�&�zp9`|�$��s4W���(ZY�����M>�԰	K���������ݓ�,;�6uG����uӫ�Kg��#�$A��ͬ���hH�p=R�u]��c#��+xaY�O����n�%j�������-����T8|�a��#':6y������9�n� uŒ�Wsro���s��21�|��C����A��꺡��u7&&i���Fg튙��N'D��%�_�0���˳0\���^��uM"6rj��,�U#G�B��@���s��]0���u_�Dօx(%�fuW�������w��Iyj�9A�ME�����R6���26b6Lf��LXs9t=��St,�K��Y��Q�ة���_Zg
����H\1��&̰IY���co]��I�X��h�N΢K���n���5n�^2��.�N_�.���e��ͺ.����&o6� ��o��v�aia�fw(�\�S
��M)3c���	5	��LgԅJ�����2��:R����$9��7&��mQ���?B����uS��*R�8�߰ob�^t�ra�`�t� ����!(�nc�u4��t�uQ��g�2j&3��l]��j������wKty����Z��{8sT����fܜ�d�=WRV4-��|0B��1s��fe�֭��]��-�Ry=V����T��G ٣�^�a�2�Ll����n?X˿�e���0k�t��_�ۛ��2����}�AJ����t�;��ȉX���a�f6�YM8ҟsw��ٻL.�J�7*���Tx���`�{�'�:Bݩ}h8�/�~bV��f8(��.�q����1\�*��Yr8�V��^���L���>����~yuy��s�����ro�,Y�)csz�Yg2�0q,^~+w1�[n�yÀa����cp �Lĺ���q�2h��	W�c�����x���wa8pǐ(J�5+��&fҿ(u�խ�|[
1Zr`	.�n���.�o��IB��.(��5\75f"֥B<�,17�LԺ����p���<�� vBnv�u�8!�(A� ��I� �07_̀0����O�#�˪�f.����jV��jt3`
Z�pAs� sJmn�S���m��Ug؃&�y�Y�,b0��;SVr����&�Z4j���EsX6�&ja�ssh�D6+7��)��#��U�Gf}ڑc�<sYp��u�6<0�uK��ff�e��#fY.�n�sn�.��d![�������l�LM��%񚎲��'���3���=���fs�D�Hu��:/�e$'\�Ո���yuFǩ�مE̒Y8-���f�N���Ó���=WsjF�+>��h��(�'�e�n���8 G�3����d�������B�nU/�8'8I�L�Cι����0y8�GC�H�Y*�e����⟘�~�#�+�=S7��/���Q��o�7���p�m�:�o�>4b�bF�hℷz��cT�E�ˈ|6���e��bؘ9Pˠ�ߜ����fݓ�[��[r��T�֜��2Tp���F�v`�$���^m��lG&���}�9��4�6�X7��2N��B3����D����a��.4��Q8�"r��mό"�"N�@mJ*H�<a�dA��X_.`�%WsQ�9�C���sa�!�0�fvW�L,f�m^�Q��Ĩ���彶��L�Rc�:-�ٶ{�6�fcK�Mr& 9�TΓW�n����F�$Z�%��e gCfڿQ�ꝟ���us�7�.6n�?�e��b^r4a������ݸ9�d�4dȰ3k&g�Vf�m��W �1Zݽs�������:7d���n� 0M��Df%V�t���c=6� p��f;�8��)�&�M\dh�W��p��+6�$}�kf��࿶�S�f����KZ��rN�n�i7G�=s���O��҄��K�~v�<�} S�fn���=7I�"��35��br�~1��9N�,z0'E[��]�6��51�4�� fc~�6���f��$��pG)7h"�ҭ���u�4���sٟp�:9[�Y���Q�&��se�s��Y�ͱ�k�@sF�IZ��^r��q#f�u`�T5C�s>�~�X륵)3lF�8��^2Cs9rk��[(�N�$���ͻ9 g�.\�$f�YI71h���/&b]�t ]��`��w��&�fPT��f�(Аs9�Sx=6�h�#c�M
���1��Ҏ�'3�:b�YX�t�	(�zf81ƻ98���6f&ZY�UB� np���	Kj1G�&o�:��.�j=O2��bΘ���A�ɼ���s�����2�"S�ܬ?���9y�İvY�s4pT0Q벬+��nx�N�0�?)�[5pؠӬ���=�,�$���-<l�li���$��R7�G�P^@h��s.�Y�����^4�m�FNL�=>���.��u����L�����j�*8���vr��p6�yV6�N'D��%�_�0�r#���ˁ�0��aE9�g��徻�K�L4S/��|L��H��[���F�vG]���+}� s����1@��r�h�9��6�n��Up�2���-d�e3j"�04g&�UV#���7sD�q�F͡c�ՁSa��.k�<ǧ�Y7�J4�f1��xa�,#fY/�nVu�����G̚/�)��.�5\��m#dj���a���(�Z���h0獙aD.��t���5B��L�v+"��-<1��@gɜMl���QΦ��Qs�aӅ�/���u^G11�[��}�Ԝ�Q���8�GY.�d��)ƥ�xn#W;� ��v�볆I�,��]�bܜuSx([73pNh2p�x����i��B3���@o4�/ۅhq ֶa����fN,7n2�-Z7S.���zE*<^Wq�ަ��Y��^����\}]o9�b��h�0.� "f�D#fy���G(�pŸl�#c���Z-:7�>k�f57r����<�m��	W�
�������e��#�̡��m�Lx���8@�9q�Tx�3���o��q������������Y&h4\"�c9x��1��M�L'D��%�_�0��4 M����G��_�b��9�ʩ=�2�8�{w����+������)2���d��u��E�*ۈ�[;4!S7'0�uE
|]\�G�n�:�CF�C� �����7�P5�8-�mN�d����v�Ո	�¨�G�1�e�KΞ��fXT�P(&,�Q-�(��!�+gd�FN�pAG�E�i3l؄!F�b�i���vlܘH��e�܈*����M��*�	[�6r^�Nfܨ��M,�5\~[2j2���_O8ۭ�4S�
k�f1���'��m��(b�:��+�t�,�e�]¿Ud� �E΃v�2d�F`�&s'�$�/�r�%���܅��Բ^�� f�����0��
/�m�$��PGf�����םLҺq���2p�n���Fǟ9n�ƃĜNd�D,+���U@s;>�	Sr5S�� *L�m�9�l��qBS�)5���7U�M�$0k��Z���¶�n:����3��I&�n���Xnp�|��H����� A�{�f����5e��XXFl�Ĕ�9{��!8�)[�-���1�nr�'�i�T�rd��q���MXRݨ����w΂$'Y�J?�ù�l���_>#�S�1'�:�q3�I���Jx�(M�_>d��>6m��qW�^N,A�	l4`�Th�
5��J�-`V�͡����s�-�61�Z��� ����,�k��K�lc�4~M�ܯ�u��]xȐ1���Nҿ|,���t��qBj;P�PA��	���f�0\N��dq�q3Pg<��53�ζ�b����p3��YLK�>B���7IH8"ќ���n2!R�f�{~0�1(�q��7f}���F� ��X��c&�kݗ6����mn��!P��h��@��f�B���['&uQ��V�>�p���[$�[Pkh�[9o��>
À	9�ģ~�6�ɫEk5n��9�ɸY%6�+�A�ZG3n�t������FɀI��5\JK}�7���4�t	�y�d�.�u{�IX�,
7l�,8r�K�z�V�-�����+��`6C�N�Iĸ���[�f�N-\�e����
��¥�t.�r�FM��(�p���v�d��3l��[��S/�G9���&����[]2Q늟�{��ܮ�f�A��Y�@�s�^�E�@����M��h֎�2.j/��ɀY��I�a�uY��M�q�z��t!C���6s�->�����+�0	��K7�x��ήs��u$S���:��l��f��s0莑f�`��՞�hu)����gm܄'�a؍�Q�̯⾙��퀳��I��9lΟ�Ϧ�k=b��S����Ϟ!Fh�jF9筘�=��)�𑩰}��+%'�h�Z�hЀS����e�{�lDL��Y�p��u�d_�d#�5��[&���`�,��A欈��a��Z��́w�/�Ձ����0t�
�}
qBj;P�PA��	�, ��`�����Z,�����Ԟ5s�KWP f&�pō���Z�)���ѐ9�ց�B�]� _y�/H9n�T�����o���)��Y#5/�'g�<�	�$�ט�5���W��V�hV:���*.����]L��"�z,��y�^l&\1�,��'7gA)\����l���2�9���h���Z�n���A����Ԝj�Y�5Q3l[��$To��v���6d
jV�z��ԙ���-�3�]N��/��F��AQj����{��,o0p�f^���l����1N2rnyUy�	gM��C\�!e�s��ɠ!�&�[��e�6�bi����j��hЬ_�ͩY�5^�j��d��a���{=�t�Q��#�$H�?R��Ǜ���\�2���+� }�b<��V��"�B}��l�Wq�M�K쾩QsB�aS}s��L|4g��3fmfy-Ҥ3
/�p�4�͆�1�\��r��B7��!�!�����6��7�2�6z�X�+�*�����b����?|�ñ�}�]���p��)��뾰.��f]P�������L&��8�ٜ(1���=��1s����e��,pj6��bj��kp/��$/��9���w'ja��9p��!�#�!��?+��tuŬ.�����8ou��$J8#��r(NZ�<W��Y�b�dR/�W���ԌNnԬú�Y17l�f�V�7���pň�����$6rؘ�u�8!�(A� ��I֦� ���z_��<UO��s�/��f�bf���m#�X ���m7����p�=	���>p�P��ef�uq"��Zvn��`s��I֭�0C��"#��ɑÆ��ͬ�6j�|/\`Ո���M��
�d��8�$�mtu��ㆮ�2�S�L�I`&�ZĺSu�Mw��#ǅ�۹6˛M-$s��n&��g�W��9�������ՈI�n�ܥc���
tY:`�`0jnU#5t�PV�y4hԬ��/!R���mV#�,K�C�M��fVy�h�D���̺�a3��D��N�b���*3��bQ/o3n��	=Ĝ�r���-��p�F������ˁ̦�s��fУ�E�p�W��a栄FN�+P�-�`��ۦ�s%m�HT�K`�j�Mĺ����,26g��/<��,0rܸ9�._�3s9K�4�N�p�ǧ�Y7���t<r̠q�&Y(F̹��h��)���'�vk��e%��Ӵ����u_�� Lc)�fA|�y���TuH��:U�$}�Tx�݈9D/9a���y����>fbT���C����2_�Su�uL�,9<�5�~����9~P�����0Ÿ���3ru��za����a�-K|��^7g�
��i�f�	MN��~N��oV��tV��$/��|�kv���!c`�����9̜Xn�d�[����ȁ��H��ٓ.���4k�ޫ'斨���`�#�8��ƃ�"��>�l��x��	W1����lJ4r����:ĀϚ���F.�����܆���p�Y�C5�E��'y��;��m�db��`|�\���h���亾�ǩ�f�,�KBL���+6�|��y�pE�Ď�R�FǨ6E2E���� T�~y�$���0\��9r���@�C���sA�!�БYE3��jfB��"���Ȝ�n̘���,�ܝ�P�իsɟ��T����s��$���CԢ��PSak����̓�I"�
P���jlv�Y��1[�D�r�3h�D-,�^����Q�M�bl�!fm������	9��g���i�9h��Z8ٖ����$jց��} pS9"Čw�����.��(�?@�79p��MI��so��S���|�qs�@�6���]P�)9Q��ހ�zIШ�<�ㅧ����S��f��,���jn:L���j�/�ب���J.ӥL&�W5�u�Զ�Μ�d�%8�<2I�?���;����V�V.���3#�294����Q�0e�6�|�Oi=�Y0���DXåd�n�<\58�l�ZUGܜ�p��&��a*\�{�,ߥ�t$R�1r�,�u;+�$��p�6�.;07wm�;���l����F��uh�b���R��#Z�s��PQ��{mk���V��E,Q� 3X��O�L͕F3��5u�<Ĝ�;%�%:،�c8��N����r���%��܆S�\�erGV�	��Z���pl|5؈��0���-j.��/P��G�Q�摊#+���E��M���
��3�t�M��,Bݪm�,0D�j�KAΒ}�B��p4���8([�˟̕p����Z���<��#� �&L1"��9�gÆ����BE���� T�~y�$�*]~��r��Y���Pʁs0�S{V�
&�1333��6���G��r
0�g9b��'6�����\�s�Jl�W���W��Z }�G�EX�bJ����^ �$8t�_�ON�������M#��8�]�e��Q|]6��&�<p)��BtH s��$bl��\|��PR��l6��KF�q��s��eZaۤ����\�O�d��3l��[�Q]��Y��,Df䤨�^`F31G:2Q늟�{�d>�	W5S�>V0��nB,�5���M��֯���c̢�M
��Y�æ7%��5�<ٜh`bh��Cs���Z���	�|&A�{�f�u9����+�H&��%t:���:1�9�����iO(0��.��z�������?Kܨ���*�fϜC�9��U>Ο�Ϧ�f��p��p%�\*6n�	G��<��)G����d��G�r
/ѪϺ�9CN,>�ll�V����>���^i4bb��J�ʅo���̂~1�y��.F�k��b�,���e�DWni�1�<,�(+��P��~���`���s�.��jf醡P'D��%�_�0�Z^hv� ��d</�2�JN�Yc0gϱtլ��z=�p�t7��z��9ݎ+1fR���z�Yd�+�����z-����$�ˇ�Ն3�W��Y�jɡ9Q��/\nr���y�3j����}7	Y_x�ؐ��z��S赆�t�( ���uϹ�븺
�Oȳ�3l���=KnC�������/%5Cm4	V/7.��Ɩ]���z�����D���z�W�fЄ�P�:=�\���� Z�f�$�֣���V_͕]A�vuS��}�e�i����:�v���H��V	bBj������hn�:��b�s�e�"�my�E�s�\f�c��&d
�p/�E�%Y�n��Ѱ�d�Ժ��as�n����,�.���ͩ��%�:,l�?��:�Y.��F��97k!�1y�a��3R�
t���n�$Y���� �pUѬ��#�4XgG�tE�n�Ժ�y�?o�0�Iԭ���̒_�n�D�U�<`���\҅w;3oj���~��S�"�.ȇ3�
���pp^.4`��\we�sq��h�C�u���`�d^�����9��p�ԺE�4X�Շ�7��H��yw�r}���MJ�.7�k��9K3+�>7��ڥ��p���+�,(1�`f��Y{0lR ��ͤ�S|�o�S��d�H�7oe7m�-�qH_	1G��c&F��d)ȹ�n�0���H���#C�w����r%#&ja�ᱴ2����0�8����s?�TgЌʫ���O�ea��.�6fj�0�q8o2p�x^&��e��A�h�E8K��H�9��6s�.70�����с:��R��PI@�T��h��K��?�ݠ��b�@��]�5Z\q0���,'2Y �>��7�S��e�`���ݙ�VgN,5G�&f�8`�ŝidf��֙��څ�p��L�1���$y��HX��鑂���� ����p���Ϳ5F���y���.�p�h����Qذ�N����gr�J'D��%�_�0�b�m}��r\��+�]���ԞYXWrw阹@�bB�9J6k�,�ՒS`I�A�H<�S��p|�\�Ub��m�j�C��5�[]�j��/���g�7S��+�����d��R��C����y#栳�6)b���@���`S
�T�lf�%���j�9�����2]�C����.�C�	f5I_#.ȫ���ׁL��q���p2�~Wp�wcFN���f4#f������W�BY�[�	W5S�f)^ ���xNC3�>F�j6��́i_�^Tl��mw��W3=ǰ��qSb�9��'�Lm��5;D-���忉j�>L�6���:�r*bW�+�H&��%t:�+pxV��}$#�xB���hu)�7��۳6n�0|1�<5��
L�!�d�m��������z/�c�d�7C��#�
7��E����d��G�r
�aS�Y�k�!'�h�o�f��U�?��J�e`V����LU��_2W��^�a��ʋ�^.�璜�[�gE>�'ʊ�9���A��v�y����]�����C�"N�@mJ*H�<a�D���.'�y�X��@�Vrj��9{��+�j35�3b�uD��jh2j� 0K���a�p�\�C�For-ܜ��8X���+��tثT_h���Ih��G��s�,!G�[�+�&&B��M�h����q$R�!T�:ݖŞ��RX.`V��꯿������M���g����gyx`�y��+�:KFL8 ��j! #g`^��p�_w8o�So���nn�/�տ�`Ą��;lnR!G�[e6��fSk��L"��q���|��9��Ѻ��q#'i��3�`�.��`On�<M!��C�J�YY2r�	1�W4dܸ9���R�խ=�vc���f�.��GN�3㫙��G-���;�$��V7+�i0`l�W�&�9�U�(�9ѯ���Ь�e��T���[�u��1ur�'6d�VΆ��[����ڨ��2��X��8��L���#`Vb����*ra��Uv���_���81ͤB����-�l*l�q�\�u�������8A�$�,R��]��͢��unt��Y���H�v�6��u\Ť��!s�]�%V�Z�������p��G*�s�̜��M� �*�����FL�����ܺ�I�4�\�=2`�9f�f_Ũ��1p��%��H�:/��6ٙ#cuh5k��{�����MJ#��2��o&F/17��uh�S�94�U΂%F�41z�a�w)��!#'ja�k�6�)8`��)҅!F$^.�nv͜xh��.�cu�o���Z,n�i�$Z��Mɹ���$�����2F�c1+�zo����/sG�&���L��9$�	K�������^Rf�#�6�����	W��y3�?8�Q�dj��u�6��e'�p;s��(��/ΐ���ܨ1s�W]NS֋ڍ2��
L=���#���x8@sq��|*��v�����&Y@и��X0�ay�9���Y8p��S{N����^% fj����?�&ٌ�j�,E8�q3KZ���Y�5_m9G41��I����|��13k����h2]�~4�BnJ5���pcf	/8��U\�K|ĢQ�$�
Z�`�,�mܐ�ZW�4c�m#�<0�&L�쎴uQS!l��漕�P�B8߳n`bX�N�*.���c&���4`� 6��>���"�l�fVr��ú�ڪ��+��J�w3I_�t�W�̼7rj!�A�Rb�N�N�m��,0'W)<a7��4|q�b7�^ǆ9ř����c�ؐI!�hN�u8l�T���f �CAX
�ꇜ�*@d_#�Y�ܬ���8?����*F��.[����9f�$�Ռ��y��nj�]4b��yf�,�$��9�v'2n��ɰ��%�WM��C͒Y��K��+����<���$Wq#b��-S8U��u=/9rb"��Wl5�uh�򠼐ɹ\1���W̩��Ȑ!g�E^�hc�n����=|'U��j��́�M�pT-�[�vb��B�|�g5w6�f�A��v��f�ęv=�qS辉5�}��T9Z�=�����eǀ�+��3�M��Ε^��=�Z�n��J���P���ϗ��ȅY�Ky�^�%�&l�ޥ��lVNq䤅s��jb"���ƫ���t�b=�����Dƌ�d����6�����f�{~��I_Uf�O��%ja���U_rd�q
��� ��qo�d��Y�I�D+\�`��B�FL;"�9����/nbر��r#��b�ά�1b���l�,f+!NĺT*8d��b9Q�r���P��pSx��Ž��qBj;P�PA��	�, f��>�p9�͒=|�Y�ZN�Ynƭ�\������ |*�h�Tj��C�ٶ�I�#.�U�E3�JBācM�lr�v���/1bШIbo��&9o��h���`�j�/�E��&,1^x$lk��KL-�`N1'�rM.�E}����.�u:,��0n�p��7�t)`��Kkc��f�SB�n�`�՛N¢�f��v�,6	k���4��M
��[nrb��RxOŜ��N��0�`��B�x�o�&�ӑ�4h�l��p�0-j9�I.|`NA2���ň�ZXh��=詼>�:L1��23#��p��!E�bܼƍ�!<3��E�8�6�]N�ׁ8jV�S->��Ez]�$#DC�������
3�Z3���̊���w��ݒ�:��ύ��g��M�ㅛ_׃��ǌ�Z��-�}3�|G��͘Y�S�?Ba����%�Y��1&��ɏ�mK5+���s�R�_g��n�dڀs�.h67=�H�W�Fϲ_'4)#�:�;D�
�I��-ެ7k�f��"�_�Vf�hF���ʪY4b��e��l�:�A�7�J���̐Y~h�UN�J'D��%�_�0�r$������a��3df#��<Ҫ-dV��=b��>�G���fS�����m7��/f�W[��FL-\R�5[ �$D��f�fg�!���"b�6k�'<��M�h�T_�>�O�u�T�Wك��$�qC&j]�ӌ�붍2��M�"�9�o뢆��b��}���"��S�¥��R�������
��#M��1㚞n��15hjᚳ�s�O�D���cf��W��u��J�9��:���<3R7�w��|�N�?��4!J�9�|̬�K�XA�t��)Z�3���i�&F�cP�ax	_�.ds;�Ir�M�:j�=}��Rf��TxXsL,�}1b�16�̾a˭ֹ�f�^t��uf6��������;3�x�I�����l�D-�a`r���ȅ%��+|Ř)�n�fm6���$3Ռ�nVtݖie�b]�屲�OM��s_�K������9���Lf4ƙ@���!��9�5q/�K�f0X��|��P4������pU�Mq�)؍-˵K�d��X�s��Z�1����^��S����'Œ\ �G��"a3�I
=R��y�xԛI�j�B4`��[�bذ.p�,�����ljẫy�ksb��tp:��Ռ\��~~l��o�"�KF�6���4W�z�!'&¡��:�w�?5C�u�d�d�B~m�������)��d+���̾��S'ja�����q2��p�8�^tXZ��.Dsq��$�ṡ�p�Y6��vIvD*T3��h�,�`bر:�R\�K�Lu���'2h�$�����_)1p����y�:�9�#�����"�:��p��"��y�.T�	��@	B�'L�6�Z� ����Ӓ ��~<�L�Y��3í53z�r���4�v�>t�b�к$(�p�'�7�#'�Vg�"�E4/�P�|ѠYh���,Y(纻9�֡p�}�]��Ő���.~1l�����^(�z?$<k�p�n�6�/Ӛ.C2I_#�qGα��ΘI�rݖ��t�>ˍ�L�+��p#M�W0/;nM���G7AL`�B6�f#�p���Ч��E�r]N�����^�r� �L��X�o�F�$
�e×��7���4�JΗD�=�m�l,t:ϖ&�M,96j��/\���$#󰅵fN�gg�FNJ�nf��\�s��i�%t�O6I?������2%3��(�J7�΃��n�p����I���6�q1�bS �49�x��d1kjf��Yh�D�U��M�����tȜ�#L��s����s�	_�Qxl�9�T*�Ya�+p�<�$9�����%{��p-��EW�H�y�i�s��y:���[�%|s�t6��bJ��Xc0lԐ�S)����s�nks�u�fY���s'Lu��2s�%}�P����םL��;p^,6nN�Z��{b^��L�Ĭ�C�ݺ�a�&ja�̲�^79�<L1�H6bĀƫ)�v��+�&N�f+��\7S d���9+�nR�fV�>�Ny5Em8o9ʗ�Z���6��͡�8���硋�!%����j��2/f�٬��LL!�Ô�!���&"l�R-��[�'�����e+��s��/<���3v	�\ѥ��Ň��H�y�Er�ը)���f���U�I�G+��r[�AC��#�
�6ǔ�c$�i`�c0��+�W�-��>�+�F#�rQSa�����w�$1I���Y.+YxtwO�S�,c#d2��\<�U���ޢ9͏��nd����-܈YΚ��p�~nr����c�q�BE���� T�~y�$kyl�`Vc]��%���!���ڳƇ/2�fv� 1S,g��Pʹ�d��'
�#���~����MQf�cf�i�C�p=�,��[4_�u�q�ùj�ȩul�����a�d�����X�uvS",+0+�0�a�&����:���%7�7qt��f�$��T���G�;��Lґ�8n�-�M���O9��LZ�<�U�5�nW��ѭ&	�h��Hr�6��輊B��(��nKra$3hSdcc��F������-�3�.�p�]47T��$��YW57b�����Y��uf���|9�l�ZK�M�7�R���$'��9���q&Jẟ?�T�݊q�v����<������[�,}4Ip�b�o(5���|u�4-�s����^�dVz4l�Ɩݮ��b����:��s	ov�
�-1�fтI��nA1�f�7��sap�:r�+�"d5�9B��O��'�J��긩�~���Oa4I0�,�E��	1�O7�����d�-=�v�Y�r6���-8،�k����Ff���~$��Tgf!!��2[�	ʍ#��M/3�p��1�F́EL�NC63b!p�t�
��0y��hL�>a���m����!w3b�N���u���rh��Y�]0M�ȅ���m}�����pg�ྙT�/\w9j���/�jj�k��h��ѕ�8Z����,0h�$A1J�u�^�E*'�W3��PVSh�^G犩̺ٞ�j�Q�f���;`
�pn�"��ڑ
�\�u�sxL@��,�`�1n)\d~�lNJ���Q}�c�LF}|a��:.�h��̑��9�Hn2�nd�9P�!��3gA^G2�᤯Q
�,�5j6y�%co�w�Yn�6g�;6j�"�I�u�<�ՠYy2Q��덦�E.;��V��ڴ�$S����%G͓U�L�Q��4I)R����A#f�	'����r9N`1�RO��K6�&Kn��>���Z�`��,�%�&\�l����Aj�b��5�Bp�T��/5f�\T9`�$��T��j6��H1L�s^0f6T�vٙ����^N�>�ee�<���0��M`@Ȅ+F$Ο<��B�0xS�	��@	B�'L���i@�f��p�0�8�LN�Y�����?4kQC�tÉ,����:zN�͝�	���6����p1n�$�~�cA��vx��{џg}��Q���&��5�ʊ_��E���Y?2l��%%Ǎ5{�LL�-q1'i�M�jfN��q��qS-Z�ǣ53��M��e��Y���j�3�υ~m���)yʁ���~��5�R��w�R,�����8�f��a�H��0�t�Ô^��^fd���3��M�9��~Sw��i���t�W�͵\0O��uſs�#,�E18G�ˉ�v��_� �9�mt�k��ܒ^��\���
�����sb���$�$��0�L[�rhV��|~4r�$y�b̜~f��j�i�/>R�6N�eP���s	���d"ԭ��;��܆�Y��\��ηv`��[;�G'ĥ~�?Fb�����6���d��K�́�(X�� �F�I���=��D����p�uO����P�Mx�� 9��[tb�<��;b�����@��/�������3s��;ne�z�f aɉ�X����f�]Vh0L�#����ڽ�M�{E����'L�6�J� ���,�KyH�S{.3dn2p�h����ͥ{����M�F��(Hشzr���WEM�ݎU!#���$1���l1��_�^���-^�$������UM�f�W��ڀ�$���ՒD�|���t}oٍv3�O��@�zm�̕N�~����\�`�t�f���ɺ�]��?Њ�
��-��p��Ĩ_���D8��Iќ�pF�[��"'��a�{�8%f�@	B���L�eH��̄�8F`��C���k�UdS�J�s��d��e>�S݁�R�����߲�!��,�uGs�m���26��u^��XN���z�%~���b����LgO��:41�i��{9�Y��;�&�^�FN��Yh�Trmj3��N��_A�E����Q�V}�����L�uw��7��ϭ�s��!Q�fr�y��T�F�˾�!�fy����t9�ѫ
�����uaw#�;/�̀-�U�0�P-�s�X���H�)5���e�N�6d�7Y��+x���#�ݖsh2s�:܈I����<�5^���et�ms��������nQ���)L�2/�M�Y6pࠉV���F�9����p�>���>��Tw�ͳ�PkFN���XίS��j��s z2I��]�å5+�fH�p;R��K+vlİr�P؜����p��\���K@0z����up��8GV
���Z�{Q��b�C�e�l��M_��K�Ws���.��R+!�`�Ġ���Swɵ��~<�1���
��϶��͡XL�:E����'L���i�����;�k�zb��γ�{�l	-��B���MvP�=h�<�5U37l��wF��m�j|>O��O��*���4]̺�y��c���ܩ9p$�N�E���'���ޫ��e����K��l��as�.�Ek�f�*fюx)����hSP1���ں��RL��m8pbN��#��͚.��7u��+�f�|Q/�ʸU=P薰�d�·��[��M����;��&E��̼dy���;���uU��ՔP���
�͑�aOU��ke6|~�!S��e۬����l���ک� ��+d��Z0	~�Za2���WS�>圙��I֝���!��n��-Л<�&���%�f���, |�^A�dиq����Wv�ќ	.�]n5dchR�O��w�u�|��kY��FO��R7ja�A��|�$7`�Ĕ�1bR�WN���y�<���f�a��!j2����6�d8d
��왹u˘LRX�kX����֭�bEs�\q8i��-��̗�ZһQ3���a-M6��r1f��g�����'�6zv��9T�>-���B11б����.�f�T�����n��n���u��,��L����!�Muݼno�v���g�dYo:�n7{ٲYM6jj��ſ�
�#$1g��q�Vߎ�C�Aj7��+h݆��M�;�,t�naw���uh. 6G�j�d��8��[�)��I��6(A� ��I3��c![�5]k�f���`,���}!�Ӳ���^�\\v�m~W�f�[�����{0���`��,����\ˣ��n�$�����w���(|nl���Ƿlٯ����lx�F�u2��;�?3�s��>�S�؏��"Q�tk�a2{r����p�@xR�1c��Hr���(%���^Lђ]�B�������jNa�#f]Ԍ/�P0�����C���UL��+x_���!Ӳ.�j�<�I�L&�ԉ9���#�r$B]�o���sz]8k�&<�7{�f�j�a���{io��$G6���{"/��*��:�9��I��,���妳�3�`���Ԥz���Ki�ϋ.[���T�^���n�\�M-#8���]^�WJL�����܁j7Uh�S�b��Ո���A��L��P����@1B���{�l�D��\_6k��M�R/d�rA�(0�n=Ne0o�I}����|�k8�����N��b����Ȅ'=�l�v)����k�f@�pXU9�q��1j�|[4b�Vc��e��p�,�e�͊�	S��Mr0��n�d~�Y��h��G�S�	��@	B�'L���Y1}���L3�>|XP7��4ݪ��YVd����)�?��9��,�-�LK����9	ۣ�=ݪm̀u�G̍�����(_�%�&3l��ߨ���rj̄'�f���J�)�3sr_�7����UTs����N�:7f���{�D�͡�ח��A�Y�f(B���L�n���fCh��!o�n�I�4?T/�=9h�D�+�_#2��/�M�ҫ9�������>�m���Q���D�#V��!f��q3$-���Y�lf��T��I�N)5I���=� 7������!3V���:��,����,:$]�����
-z�ã�����.Ue99�]΁��w��������3I�E��
�aY_531GsW߅f��uͅv�s�����p���%ˆ��u���Af�n��	S�(|_�ۯ��S�qBj;P�PA��	�, +d�0�G]0���$��h7-8f��2>k�w���>�.�M�+P�y�Ŷ�\=9	�����g<��TF��nY.�f���M�X׆mt��c��7��ԭ�m��GMʲ���붗�j��qvV��ɺ�#�,�s��tݚ/�t&m$Lu+�xD��������l�(��ޑI&_PϚ���m�u\�98+�&��Ͳ�3f��
W7�y̰Y�p���}9?�:-�p�THZ�Ml�X���ο���W�X�m7q?��P��#p,B��t�����Eͺ.�%�A6j*���fыIu��������4He��㐲�,�(Luj�}`��*m��x��i�.�Sml���,��$gxC��Lf}լ��b��0�-n�A6���>G�[�j��ѧf'����ຶ�ND�s��[��8� $E��: B�'L���9�樀|�/���Z�9���������Rb��t��,���]�f��=���7��M�i�E%H4���E1�L(���]8dh=�T�8Р!�l�&2	עԉY��vV�Y;5Iۗ�ub�<�39jB�n7d��ؕH��1��ܬ��Թ9 ���d�9]�h�,�u�#� <uh�׌��/qJ�[w��,lk���e�p7b���Y�mɄ'��������\�<˺��5C&Y��3��j�;=�I8\P��)�F�;/����O��n�����z�u��{`��:���fs��M� N�joXj� W˾А�Mäz��5b�jh����?��rs��h-��	��u%�*��nE�LxR�Y���2��b�T���� �Y^p��I�m�D^�6�E5zM�E���l0&}��f3D�O�a.��+'I�'��T��:w�}#��K��VI����3�]����uG�u#�ҙ}pY���r�@�95��MV6�p�ۦo]ĺ�_4f��u�Z���As�.�}8�p5��5\�%s��RGf���c���$�F�[ Vf�/@h}��9hVq���G s���J%9��2���#&b]��s�=�9<����b i=;fĬ��9���)[��sc�MSy�cy�_�s�Mҷ(ul��,��G��)��v�����&Y@�1}���8r73nN��c3jJ��}z%�qG��|ŏ�F�K^����77h�ZG�{�U����$#�@��,p�s�&<�r��Y5j8a0C 8ʃCX@�9��UP�@�9=���}��ѻRG�#sլ�b�d�"ֹ13e`ܘI2�u癘{�fq�i��M��!��^�d�!��	L�m{�`Z�$�ܶ3y��̪XW�[�O��E�0�_�M-R7Kh���y�q� r���nn�K�!�[�!i�o�,�+�h�T��AsR���11�~��Ϳl!s3P�4^�Psy-)3b��Koi���nԸI9�����&����e��Y^��F�K^���^�|V֯02f�����a�s������c&�_�����y)�-A�q�����M�{!�fbN�8������i�.O�ӞDl��9aJ��ϸN�G3��Z��"Pہ�
�/O�d�3��fQ�s�3�;JՔ��x�2#�]_4@�����o��V�2��Ǆ�c�CȂ���g]Q4nB��@�L�ܸ@LJ�h��։	Kݺ�yT6kw%��_��^��x�0�YJ�h�E���/3nB�oh��Ya`��@��D/[/4�!4dRѣթ1s~mέ��i�u�sr-7lԄ�L��p�-Փ�M�:1�n]�|2�$[k5��<F���D��"�͂��(��.M8K�Z����;��u��I���]�ͭ7	л�b6͕��ܛ��.fȬ��d�����J�L�^8�.fA��B�ʛ�3^w�ك���\91�7v0T���j��-�Ͳ9��I	�:5w|w�`ȠQS���^LR�e��X�r�O���[��8���$�66��'f�9�fs�揣N�Z�vQ�9��HSqR4��31��9C�� S|[�S�͝:˓�ecF�
6��k������o����i&<u��T.85�L��P{�׌�"c��C�M�!s��l�\�`.��'a�y?v<��"�5X�F���(�|��{C�������)4pb�^�G�����&ZYN����7j�L��Ū#&u�X�͉9��u�g3f�T�*G��p"�e�Wi���t��̸�fo��$����}�{�Z��ȼj�r܈I�@�"Zy7d6�̚�lV�%_�SC&Q��y1�t�$I�ni-�����ؘ��� %��è�$�Đ�����`N81����Hu�8!�(A� ��I4@�����s��Y�z��Ք�3��3sY7 f����G�:�K�49�kS�گ]���ZJlؐ���(z�l�l��ůhuQ�za�Z/9�,7j�tp3�!�����B����2�Q�"du+�ќ��������e��&Y�DYX�
��lEذ9l�`��)[�r�,+6 �����E56�o�/;�V|Y��IQM��:1ᨋnU�:6h��Brz�I�0Y6��a&���$�57m��8j£92�k��3l�U�P���N嗚�88�9!�L��Z��68���6̍��$s��i��e�̕_hVE��.[�]6l䬨5)h]��f!k�Zl9���lt��q�H��j֐ͱ�u���W��C�L���n��zt&��R7.��Scf��I�gs	�����U`�4G��8�n�
\H�����u
�9���
d��_a0������&��y�ڂQSgYnlEݰ��l�ʗ�
2��S���2)��'G_4p�u�b�E���+Vݾ�df�M�I���o��ަn�]߻-���w�}���R�(���u�������_+�\ݘ�X�9���v�4�����dn��W�����Bz�'�bK֭���9?�i�Nw4>1G{x��Ӏ�J�9�.G)ssa�u4�1��Y��r������	�yI�$�]^�X�r9+�/L�̓�Cƌ��7s�{*����']y9�c�Ѷ��QGN��8�\��u��� �-��X8���̂z�Vd�3�Kn��W�N'D��%�_�0��V˳0\��$�h���p�tY��E���u�Wb-K�u^�9UtCf�W�R݊�[��g=ΏA����h�e���,(p��	9�\�7`~���ӵ�7�ҋ4L�/�S��A L�%���
d���H�Ͼ3�LE&�G^(6�y01u�.̩x�GS�'s&n��ʙI����8�ob*P��:-�+�5I��LͲ8N����\3�O�$��ԝ���'�2O�%�o��&9bbT{^6`�쟀Sws�d��93����n�Ah"�ߖ9g1�]5��ѓ�a����b��i�n��s�q��4�x	,�5>�T�s/�����h�c��7�]�B��A~p��;�ِ���/k3r�u��b��1k��N:7n�����4Gb�����V�3��e�Ձ�(�C���㎜�u1KmѹY�j�~1aJ�lRΙ�K��_��7ɺ�t�H��un��C��>A1���xm�b��G�c���m����d��6뎦!u�<���5=�bT[�� �몹�X�}[V빑�q�-r��b�f$�]6n�܊8!�(A� ��I3o�0`�W�0pW��h�i a��5bί�cfB���`K�͂s��ܭM��Z/���,���63O��9�s�՜�����p�vs�����25������\��ȡ;Y����9h�6���M\�ͬ��{#�$}C撻Y�ǂ��[?3'��JM����p�,�a�]�����;3I�"ՙ��j�	�"�-�ͯ���u@9�]xs�mb=�3�)�u�� /���0*'b]6�?�k
f%�	S�a�z.S2��#�h/�[F&�٩3s���)��K��׳I���[�VCLQ������z�9	�\�uݮ���lf���I��jlt%7��?�МN���\�������1m�E^%4�'K��C��J�zḻ́sF���D�X��G�v7z��Vu��,Dh��I��B�b��Ym6]w,�V�$��w���ȹ�G�
aC&�~����8#Ԥzwoy��Iη��Ɔ�1u��X�����
���usq�h_�`�ǚ�S���l	��FVo?̖ƢVs�YG3͹!���y31����_dr�\�
h�a��a�����spBs
�c&z�"N�@mJ*H�<a�dy��0���,1�͍�C�6mj�<5?��
�L���n�_����M�I"�5p�h��g��X�]�&Y�@#�S���[�p>�+�YuQ�VE98!������sD�L̀�Z���t�wj*K�͙���2�NLX�6gfY�l��/�u�ſ0nECQ��u��a��sxlG����f]἟M�Աs�s4��ɺ5ts�X͵�$_��Z�U4� ��� 24fȬ��%����M�o-�rn����E�����#&b]�or��ltɘ	S��9<�A��+^�/�p�%,u��3��ئ&�_���G�����(���(#�bw�f.E�#�-�K��n�t7I�.�@��YH�t�uX��d�PM�j�o4n�M3�ʲ?hV��,����jNy3l.�e�T$s��^W5�?LudV|eʅ~i��!A|]�>��+�Pnv6�N�14b��r�3�O��"�I��Y�d܄�����`��&�
�s��#:)���l�z+�W�p=�#5�m�\�ͱ��e�If��ƷY78I>mt)����1�r����*��R|[xһf��-�j�Z-�Â�/�d�����z�� �E��$(��{(8�M���*�a�|Ši�ͩ���:�jꥳnK�8\$�n��OQ�˙8'�31V�qsl��C�s�5S�F`԰����z�;Q�G�KY{ăY�g�7�Iof}Ŭ��6p)��L��	~)b�Ԝ�d���[V���Ig&��Q��5�Z�h������F�aeI~�����\n�l���N�aPM��
\��#c�MԺ�N��sa�9��)��pp#��i��A3ɺx0s|��B���^�`�,�]F+PL��M.���v�Vq���`&��a��c�i/�ku�F�=6bb�R��3� zvݒx���YX��]��-��u) ,��oz!܊Lx�_^3� ̢<C��7�pv"�I���j[b/�j��f3�ij7ln�9�mt�qBj;P�PA��	�, G��>�py��;�z�W��D��M�)ΔC�� 1SC��2^��yKFNug���:WBM�^1]r�[�l��ҡ��$wם��?੦����=�%an�df�A1��[��9�̰I�y����ِ��ͷ/��%JBy�P�Q���T�Z����~��&�l��x_�|>`��bF�s�n�&<��,|lЬ�b�������6K�M����6��Z��D��lȬ���Rp~u��i�!����s�S���fWs�0�nsn��b�ԅ��/B��|^/�p�T�^�����:��,�$r�}.��!U�_��u{1h�e���sw�p٭������3WueJ�0�-0�� �L�34"����I���l��<��ˇ��Br�&�l�Wr��FL5��qs,F11��Y}2�75��<U�+CX2k���R4�� x|��mh����[��y�.{׭��m	��Ɠ�9Gp&s#���g��r�_�𤿜�~�->9d
k�\�u��0ձ�3���L���Ь�����%�{~�y��4P�u�ĕP�KT̂�� w��T09��u:���mi�9��Y��k�#�f_=7hb8���΂��a����y7Ih9���f5��/�r��sԚY&fb�n�v��AS��,()������z��k�����>&��nù�^��7��j���}y����@C&b]j�����MEw�/'�5��Mq�����FN���>���7jJ����C��	�z��8���!��m�P���,�Mo�ronY�I�nf�恶7S��d�?K+���p��fԮ^��]WL�&+�g[3�^��/�{�&�e5dm�rU�T�������$�Rw�X��l��-L��lr=�ܢ��z���&+Ce3l��:yd�D�����Y��Q4aJ����s8X�
�G'��9�Å 2j��Y�5W�ԍ�M/%3f��qBj;P�PA��	�, �1������ݸ9,�Y��M���)�f������L�6�� ��jĈ�|c�6Kls�AM����c(}ʟ����^����b�Va^���e{Q�LrRc^�5���U\3X2�}�͐Iֹ9+���6S\���>���pܘ9�a��o㓘L&/�ᘚӕMJ�׭̺�мN�l�+rn�I!#b�=��\�0%?&��:o�FMLr6O�ͨ)TY��n^N
)?��@��e���mU7z��y�J�e��۬�����g]^u�?�WՎ�%�nj2n8]��"[��o��z�X�M�p�I֝�+�� S�#�6ȹ�lb���Ls���	)�#�]�c΢6'e�����aL8m��cd�^8�a5IY�����"t�uUneҺ������,��u	֯���#M�����,�eȆLu}.�%p@N��22h.����Y��5�'���a��/6�e7j�;�ٜ�Kr�W[��*�5X���,�ly�ǻj����z�9�%�1er�x4�>Z*?��,�����������L��[�7�F��k�T����X�S�a�V����GN�>+�$�.Ř����5���Y���:�s��X�����Q�������T���2봢d���v��F�4��OK ��C8����f�c�`뻀��d��@���æR�^�V_�	C�;��WgC���~�3�e�Ɛ`��,Z1����24���^1	��X��$�����R�P�1�,�g8hbd_�d�Ҭ�n����N�W��-��]6-�2���q,�nilb]/p5r�D�k�7
f��,3��"v���[t'����!��;���BC#�pJ'D��%�_�0���B,�0�f5@�
��p9djӦĬ֪����.M f��pN���Z��`N:9Ixfg!?�,R0r*̄�`s�u4�f��I��Y�В:�Ѵ��;$��ŕ��\�#d�ٸ�Dc暂9�ŐA�H�0,�/z(3j
�7�
d����z.��Vu���+�Ds�.���h���I�R�P!�
��2L�",��$sw�}�x��fI��sF��2 �Ha��3n�<��dE�&N3�31��Ǣ}�)�ӋY�;���ȉ1��t�\��1�j΅k ����"QL��J�y�[q�+�o���Z�s	�-xhn�
!��ĄH�
R#g�;8�����̬���^tI��W�̷�L����V&��,����!S	��烙�݁>�_�n����C��TX�l��+�u� �Ss_������"#f���֝���9Sw(_9��!T$�#�Ea��z�>���ѵas���`Vǌ6	U<AU�p,5`Vl�^v0I�-���f����y��*�����ų	1I��lj�n�v�RӴ�q��y 2n�S#�uA�qæ֭�
u�<n31u�PӚ=^Ĳl�I�fy�9X�	S��tZ����5�2^ak}̊ބ�n;6��&7�ʤQ�~J8�ӕLm]�g��8�u�==/�:Y&gD8iF�M����n�iSj���}n,21b��.�3g�����0��� �J�?�
�+loM�M������2XԏS-3�F�J���I��W��E[�]6���x�����ZM9n�T�ȨY!�##��,g��G���<����K�k�o���US�;��44��1����n�_n��5Y�aa����/'�6�_�a�f�2]9�I`��h��.�����Y��ܑ0�B�C��#�-��>m�M��a-a7�ʪ\������2q�B3I/�n��~���u)��3���}p����q���:9�/�E�i81г���ꑹjj6�@��!0n���n����l�c���iH��s��9�95���9{��v�?E���� T�~y�$�AYL`���s��`U�$\�ڴ�'$s��?`/35�4�|i��s��������:�I�=����K��jB�n=V��N�luΧ����M������;�&	�~���6��:�7�67HM��;�7!4h"�e�n�3G���&L����[�G��j��J��G����#,p+#���0}���y�Zh�UKw������H~|wpv�	8�q[�ap��Y�hn|x���0Kn�<��0�_�K��ECLM�f��@�&�@��j,���0��ep��$��!�º���"u��fx�f�&����_�KuaSs��ȼ<�hq�~b*U��aW��uC#FM2�B�g�ڮ������7q�:H�P�>�F��݈X���gs��Yy4aJ��uWso��!S�%�P��޲$�#�=���*�<`Acˢ��
Z��]^�CN�ԑ��ʧD��gs�#G61��f=̬���^��s-������C95�1f�J`��&�p�j���,��5\p�ő�#9'�3Ģsd�d6�<�Ó~�y%�C��j0��>�����T]�UC�N���D|Yt~.@h�A��[�N'D��%�_�0�bfy���Żp,7���p"�Lm�ԅv��V��gf-|��>h��E��.n3`�x�k��`ج��3�uC�&T����5��&��jS�Č��@34f�l�$f=6�̪,�`*+�ͦ7pH?P&�ȌxjF3l"�e���ƷYW8�Qӓ�"g��#�j���_�M��nq�I����Y(��Yg8a0�e����Z�%T��~���ĈI&W3>�,�0�|��-W7p�a����t9\���u9������(l*و�� ͜=᩻h؜�rV�MҿuQ�9F/�d���n�4��\��!���#`��q��RL�Ԡ���р��]���E�&51�������]��/9��0a&F~6ϊ�e���u)���!�.�JaJ�vѐ9!�T��\��l�(&���ri�.�$��PUx�`�4l�)&,��VGf�J�b�[�l������&���mt�����¹+u�Z`R�Oٺ�Y8��Yc2��r��7l���d�C�j�9?J8�6uj�-3�>��|���y 8/e#�MT���K����b6��뱌W��v�G����B��Yҷu��-F̽[�iy��qBj;P�PA��	�, �w1}�Y�`�ṷ:f��aZ�ڴ�󍌚��
Z�K�L%30pZ�u�`��3�|�y]���f}���Zr�Tf�"sJ�1�!��`�flA&Y'�53Yu6�Iφ�z���lN8a�oٯ�ڸ}
z��&�[T`�$�_գ��,39��׸�/���&,0��c|��^ �:6���.���p�p6/V��a�o]a��0�ZbB�Z��ͺ�����C�2h�W�Lµ(u�mWF��z�����%�ɓ�L&��r>�Ԩٰ��F�uj���[y>�ɠ������ gQ��5[�G�0h���=�1����up*Ȯ���U¿(ud̰�=�k��$q�Y4��jl��7�/��_�k��b�$�{�SK8n��k�fK6��á��[�����椊�����C��;|e�>���Egٲ s���&��R��f���#�p���Wt�/�M\R9���0��g�#�	�#�Ef���¿$��01zAs�� �&<���*<�s���7��ޕŸ�t���斯�Z���Q�_�M-�[�M�ԝbr�Y�ˏ�$�#�ݛ�,Z�d�$4'#f#�mOM�Ӂ~��-L���Ef����8^509��l�&�[ß�0C��<Y7 $f���]3k��}�b���Gf1��XBGg�l�ଔ��UL�@�~+6���<Ix�(����0��d�rX �����˵�q�Wl]�������:p�9#�Z뺉��np�$�s��_[	t)�j�n�u�t�YG5��B�r<�࠹��$Yf��&g��J�7�6��mC&����2l̠�k._[8f���LҷHu�ڒs҂Y�Iߢԝ\ndd����7~C�T���x2�K��ۨ�;\,xr�D���Z�W�͢s	Ȅ)���25��pWe?ܠY�'�!1�n!!���s�^y��M���f�,8˰��B�ks`ظAG'3벡�6���v�,��/0I�_���4b�^~l�9}����I�=���Cם�7x1l�L��|�Y�.r]ʱM/o0j0h����s���ʲqS�?>�,�`�ǐlOd@�tݱ�����:2��99+����Q��Wb��To)�9ߏ��Lޒ^�e��GQL�\��{�Ѡ!S!{��u_8�w�>�.C0�͜Hf��7�1`�T��Fܙ�ܐf�k�k�L`-���0�ݺV�Zz{�gm�0���ljY��:���u�8!�(A� ��I�%�<� ��`.47'ےP�f���6�:9����ɱ�%8�cnm��>��p7K/E�.p��Z;Ԑq��f�w��q����^�Ȍ�f�U� ���Ue��;��fw�I������ۓ�SA����沓Iy�:4k$g���ES��m�>;.31uk~A�Y+-�Lĺ��)
fh�j~���)�ʋp�V�/�l.�w�Ia=Z݂��,3+ ���Rw%�F�ƒK���Vw[9����/�u����-;�ج˅�FL'7sQ��)�^�KI8�Q�R���s�/��B^N���ʛi�o�7�`�$A��rd�DN���r�bC&��e�m�/ת�nҺ���A|��W̄4S���k~��#삱��f�X�ղ�z��%��1�Z��wz��"�'[�K|h�1��RCfY]C7�ݜr.�7�	�<�a)�:��Í3n�lĄ)=��Z�3n;45��\�58<��0ՙ!s�|g|�� �����I��hn�8Q%8lF�CB��5��� �.���25���[�ȗ1�OL��E��`����@˚���p��j��������:	&�~�p�PS]^��}4.ԃݜ~���,i0�`�ύ0'�2ܮ���"Pہ�
�/O�d9��̑��jܸl� 87�Lm���Qsb��ZVז�B'���܏~'�,�u:������uZ��И!�&T��Í4+��Ĕ�q��hبY���9j�<���h� n�l;5ǝ9�%�I3f���Irw�����u�&b]��./�U<�=B�ҳ�4��x�©0*���f;9jbX�����݄�h6g��n����j�b[������L>��<��2aryU�K�1p6���]=�,�%�&<�zPt�.�տ�ws޵)4I��TwU����@�n��6̒T�ڃ9=v5hB�컙�!��R|ّn�`��,�bb8r�g�|5p*5��aU��C�51����I�T�O�eY����y��l�.�7�R���O��/K�ҫy��.��BZ|KaA�uI>G�{J5�[(�-�$��P]X���Cfݐ�edF���)������,]5@���z8�f,W7f6�h�,[�5Ss%��k�
?�ԸY2j�IO+7h����}1.�%������}<iМ	aJ����̲]�p*��̺��
zC��V(�U_�ըA�&��(ua��"^846r����u�8!�(A� ��I��R0\�#�����yX�Vd�YZ:�\ f&8���,�%�7��܈��H�[��F��6��.;6y��喬k\,�G��u�� `�t��4��ߖ��sP��Mױ9����f�u+p����é�/���q��k'Qg���4��7ˊ뫲'�ʫiÒ\�q��d��֭04�������7������9_ЀI�3b�A�B�?�`0����bVr�c�ùȷ��'g�wn�c��8��6�ѨAS9�������F�9jÓ~�=��	9nj��K��Xj&ɡS�:]c9�}1���3�}8nb�Ss�օ������\`��z'i�N͚�C+��d��k?�~����/�0�b���/�u ;�~��=G�	�$Z�þ���Q�%8g���Sӯ�f�j3��&Y��������#'b]&�C�9�ь�aJ��o.u+��_xsLj7f�KKl��4b�����cRG��r�-�Mn
�2�I��W�r�L�#g��-Ū�1�c2�����Q~�Yr"�e>�Y�'�ʯ��0�w���o�J�q�B��n^�s/Y5�N'D��%�_�0�������b�<1ۢ��rԔ&9�>����Zf
z���n~����{�o����I��n�7f��ڨI���b#��#'<�s�^�uY�+KFMx@f��}��0�F��?��D�$�T�9����3t
O��͋����V�:7��s)��I�?W�`���9d7���E�Y5ͼD݂v:0�AS�N�����$���y��}]�D�+�/�u#s(Yh؄)����	��_�\�r؜�ju��P�Y�`Ȁ9��iK���P�f5p
����b�| J����h�_�∡��X��l��8B�f��13�RE����n+�fS�9����u'�����g�l`���n�.��E!�L[�Ĩ9J��U3C�s]���Ω,���N�1W?�^�^C8hV��#�e�ݬ7�b�q������2�f1�L'D��%�_�0���è`��9�-�K̶��P������
��o3f7���\ǵ+@��/[2l�aI�I�}��,�U� +��Pw��ld!�ƈum�.OgmW��r`��s�f�<���U�[_4J�v��ʴ[�5k'GL��DG3.���`7���:�Y�0խ�B��%p���-�X��b�l�pKf)Ǹ.���S�1���tt����Ec�R`sfn�l�UfƢ�2��K'&�:,����Stݚ��8l�d��9����v��\a0#���p,B��t����������ަ�sjԈIq�:3���[�f��u��&�<�T��Y^h�\���dИY�yaQ�����ByV��M�z�d���8�uk��u�Ĺ���jV�ͩ.'���Ĩ1s���$�`;\�9��D�?��y݂���)��v�����&Y@�AL���l�Vn6��4���FܘYh6�ԁ����sD?��;�L8�x�ݠ��B�2��L�u�E%T4���E1�L(��LP��庄帩@�)5h6�C&�Z��%���,��[�j��/52�t��vQ�	��%�����|���-����u;rj���l��8R$���s%ؠ���n6� �Y�M�D�07����$'b]6~�ݬ��	���_v+������g����ab�,3d�u��#g��tz2[�in�Y��#։� ��?8ۉI��N��+%fq����M�베¹���M�92p#r�Y��6��3i�Ζ�F��S#`��=�y�`\<�t2hn䃹9���#�B\�GR�������ΜGr~�k۝9b�T�ѐY��f�B#'Y�xn���X71���C�=fV�ML�e}������hA_�E���I�oy�9>�<\)�o��xXT1V�9���è����c��Ͷ[%��f6{���k�qŗ�f/$61r/h7m����D����_٥�p�1Q�r��x�/�k��M���g���&<u[�!�F� f�$HG�;�W
�2%s�����ܑ�6\�Y΃���Mr�\4+%�Ȏ���[�K�t[^rؘ	O��#��p�4�� М�xL�n�>��ʇÅ�!�s��-J�)�f����R S�qBj;P�PA��	�, �<� ����t#�b3jJ��Mo䐳7pd���W���p�-���.,lr��7h�ZG�[���
\�Qc&a�ſ<��.���Kn��'F�0��X8�,����l��A�f�ms]䨩�^7��	������������d�"ֹ�\�vf��~�
�f�'X��fԐ9T��s��!�0��F�A�0R뎢���$HmrY]�b�F�+ꭒ3��S�0������I�MM����d���$�;��b9`�,7C���&��:�y4��8��x�`�$]�P�f�G���C�尮�ꯓ���"X ���ەr��}��)��P�����9U�,�d��"����,{5f�TVo��±T7vą�n���6�F�3I�"�$��:�Y������q�@w�5E��Տ���^J��pmMFMĺ,�yw!�B̄+}<��|M���9��2E���� T�~y�$�a�0��%F̀���P��Vl��ĜG�c f*����fE7��n�M�h��l�?	:t������@�f�M��]4j�b6�&��ub�R�p�Q��1Ǜ�0����z G5�,�R4���E�1!�78����"�55\�~�.V5jN���u]_2K��WsL�鲻�"������u�mn��/�[.���	��70K��v�^�FΏe)��:�I�mb�ob	�Al��]��x#ۘI1����ss�v����,Ƀ(���8�˹]��eņ���[ץ��M�I���6��b��E�LUi3+�9h����{š��T��D��n���q}�$>u��;m�[�ͭ˭r�q41*-Hh��a3���X&�G��u�ܰ1�&<���\�æ�_�`�\�[j&ɡ�M� 3xi�' �̍p��/�d�[V`�tݙz��98�I�:�Y�N�%����S�,��ʹ�I�b,|�k�Ũ��:�,ޅ���8�W͒[^fN�F�V+w�o��`b��@wf)���������t�1�[o27�$�#'b]&41K��I�l~��c��9#K��q�@39��,gcdޣ�� b׹Y߅`�}�&�G�g��W0,��L1��/���sx;��13��ll]��|�o`���pK���u���o#���aJ��V^��9�B���c#�ڌ�Z��"Pہ�
�/O�d!�b� ���a�p��،�Ҵbf�j��O=3]bؠY�K���N������A#'a{����ͣ���$\��Abܜ��9ၬ3����Ĩ	H�Q�|��٘��Xx�o^�Yp[��S!�̖�>�9�S�^nd����V����9d]
3r�Ѭ��H��B�,cC�H_'5(�d�9�f��t��-/����L�`��0|P=P��XW�_�{+��9AÔ�����n�������9lNH5��H�3��{��%�
B��k������_��0j�G)s���As��C��tv/׃����Ѻ��.hhR���b�3aV��ww����z{8ww�usą��X's0Xj��L[�N 0�U3C�5;��8��%���Ԋ�Q�n�57hĨQ�.�T�e�\Ĝ@�I��w}�^�9j�"N�@mJ*H�<a���a�0\�����o�� 3��[����:o��l������alt� ���e��e%'a���Y�wcEѸ	Sݲ0�e`��/���u?�\2]w�~!��ըI�h}�W�f�<j=g����,{��jݮ�Z�Y9g�u���(e���ͳ��f��ˈ���АI&_�bt8瀜�it�.'�WM�����5��WH׽}%vWg����B�\\�l�ͮ;H\�@��H��鍊Y�v��~��P���9�LT:E����2�us�ܨA��ڔ9��+����[�t^q�o�L�n�аQ�i4�maS�apX�vk%'b]6~�vY�Ժ����Q�&F=0WO�ao�o�~-Vغ��ʑ	W�A�9�����?B��>Z�F57?�~��9eZq7��up��LZ8��Ax�8!u��
�/O�dY1}T�^*�����ͨ)Mr��\��l��Lh7\N[5���ۺ! ]��4l�rȸqu�	ſ�uQ�2���YAd�-��
D�[F�f�!�p-J�怴rl�H�>6�^]�	���hI�y��J���s�op��)up̜�x�Ii��^7�r. 2�ݬ�`f%UJ�΍��h�V����u�x6l�c�������KE�����{��}6f���r)�!��[�/X�kjFL��k�q�J�8b�s�.�#ZL��(u�_1�������f��ݼ�q����¾�pb���ʞr����SfY�9����o�nn��Ac�"�H_���[}R%�G�Y���5�Jz5h��%��Ñ��6wb�����/5�f�B#'Y����q{�T�-�f#p�9�'��·��`�w���z�Y�m����[<�q��������p6Y���6c�a�^S�bĸ!�F����Sꋱ�կ�/�K��D��_�՜���FMĺ��e�w�Z1Q�r��{�Z�h�Tj/���ѳ�LK�1r.� faL�t���~��Cf��k	�ol�}}�T���v��$�Κ� s�j�ʲ�����0���Lx��/�i���{t2s�}L�B!�p9 ��M��9kWzўcn���֍��oY�Y� S�qBj;P�PA��	�, dd1}�y��J̉�fI lFMi��d1�~}� 1S�/��p��l�FL#uy�b�ݠIj��|a��+gTO;�n��kJ�L� ea�f��>��	D���s)��
#��G�r��f�`�`�Of�뾆p�l:��(u뵌~8`~�!��/R��ɜb�"��k�����?������au��$����O�0vݱ��W�� =	Bd�"��/��s���O��և�}Sz3����f*���辰�����H�;�N���ᆴſ�f!]�c�L���A�B1����ܨٸ�d1�R�lV�p��6���6��n��"�4������u��7u���6b����_`�,8'�⫬^�5\���#.Lug�uZ�+e&�_���2Ws������S���4/7�8�6��b�u��1�fA��j"�e��1�l�A�\�N�������(�v�Z��"Pہ�
�/O�d�3�����b^p��h C�nZ�����b8����l�lt�m`��Q��1[�Y�uBs����;�u_0j�Y07"u�)gȰY�� �������Y�s���GN8���u[�h��,��:���V�_fĄ��,ɥ�BЀ��k�8��2Ps�L��������,�mV�����u���u�m����.�P����ȸ��@�}#�}�2^wߠF�u2�������X�����9�����a&��=s����D.+�����x�"G��f�MdذQ�uk��/�
J�z7�Y��p�=t�J��)9_Ѐi��Q�J�G��S���%�y8jNF11o���y��u�rW�J�I�8j-�h��a3���Z&�K�ٷr+���C�e�����N/^6c��$��N5rV���Y8G��e!w��۽YM׹Y���:�R���]̂pr�Yѕ��O��i[��/U6�m�W�J�����.!4����f	./3'<�*T5��{tT�`ON��Rp�����1�Y6ɺu]�k8��#'b]�1f̐9IW�M�ү�z,q3gp�[O�#�9��/gђy�"������d�uG�
>T���Kz9p��ɲ�`b�����j��� �eAf�V_M�o`���pK���u���o#�z叉0���t+/fS!��]��^�QS�qBj;P�PA��	�, ��>����:w�݀ͨ)M+f�̠�̡��3S�%��u���o�r��3dܠI�x�:8�
3I�bs�ĸ9r�ig���%s�
�Q�|���4S�M�9kn׶p*$.��09k�S���A�"0?�$��n���9$^��Ь)�c�l`�hV�96Ϛ\�d�u�<�uX���ub�n哄T��k��h̸�XW�W#go�i't��/���n���v�灉�	�&Q��[����{��%�
B��k���@�8Sh�$�Ω.�i�8�$��LlN4+7ၻu[�u]�6�$��_f�*�����*-DWa��ʹC�?B�TG�V�q�rj���$�"�-�C�殚�:i����|��i@x4g�2\���/5j"�e�3�~�-J6aJ��+tA� ܖ_-S�	��@	B�'L���A3��0#�\�m�;��d7�ҍN�y`��L�a1������ 5���,�$PoN6W��и	Sݲ0���汢�/F��Ai�<��t�b��̐Y�j�$Y�>d����H�L�ZɳH��O�=�B�nׅL�[�s�8a����0�w�lb��l�C��\ѐI&_x6���#롦Ѵ�=��Y941F/�W�х�B�Α�^Wt���wn.�UsS!I��-�H��H�������t�������¾�I&�c<Ǣ��J�(�br�݇�Nb��-��Ps���O}|� ��s��EFM%�l\�F���UW�a~ӷp]�ȉZ�uȹk+�t!���b�7qj_�����W���氹h*g\x�޿@���\N�"ԝCf�Qp�H�C�9E[7��up���]���A��8!�(A� ��I�u�G��rH9���B*GMi��Hnܜ!h6��f&�.������mݐ	��;�6�b9dܸ	��06����g&d�dɬ 3-���05ʝ[z`�$܋Rg%��Yb'��3��;O��.0pЄD�q�,Ԝwl�:Q��g��XfrJݑ�p��8���M����9�-�����T�9���Y�E�}�;lm`�V����u����`.�Ò��_*b�Vz	.�k��5\>!��[�/X��ٌ��=jn8S(�Xw`@C���b�G���z��ٸ��o_�?�y_c�ͳ�A#GΚ�ild7��'θ���s09��I���7�2�y���6��.��LL0d�۲b�娉ZXb���5[���S�U_�;�{��TG�ڠ��S��j��j����-$�8fVvCɺ�Z�U| 5��m)f=��r����]|�q�p��:^B7gl�L�Qb���EE���!s�')��=�\�u���'�uZ��n�M�����uw�&b]�ł��p�p�Y�Q�r��d�\`.�6�"��m6��3$,u�AY� p�$�D��s�Wr�������>�����Sae������R`Q�s��j�ʲ����^~dN23�I~z<�4�����)>�ǔ-r�`؜Nn�l�9f�9�&�[lݍvs�.K9+��Z��"Pہ�
�/O�dY6˳0�6�]�n�4@mFMi�s��\�[��h������q��f|�T>�b�ݠIj�nK6[���3���W7C�5%c&\��0.T�G�ڻ	�W���.�N&L1����as��lu�0�ɥ
g�I�G���h^���N��nկ�{������z\,Y1h��Kl��a{��$��������ubڬ[xD$A����x��Yr�D�+��21�&1aJo��9�ݼ�L%����9I��D�C��C��nH^�[�j�U�Lf
%:4'���&�z�28���f1I�:��u���n/�g��n�;���B���#cNĺL����\1UX�Ӌ9W��O2���t���S�
\!�c宔���N+8�B�U�I����j�ܡ�W�Zmv�����[$�j"�e�1��As��>��^�~1�L'D��%�_�0�g�0�E��.�m�7��`7-�����Y��A��f�����r��fYT�&����%&ۼ�p�8K{���B�N4hԘC�AM�.��ub�םZ���6��ÿ��;��d�U���$���0
�̸	9>.�nV���,�.g3Kg=뾬АI��N�ʐ9�-��u��[@�,��<�儧N��?Э�9f�D�S�Ĩ�<#���P�21�u*�u���}��@�9lR��X���^�g���G��
`V�B�vI�7�`�!3�X�S�*d6�gl,YF�@�̀���n+l�<���Qi�꺲3vvݪ.���y '&�&Wg�,��uKԌ6���)�'����z=��:77gi<��J{����.�����$ i�[95Fq]͚]���1F�k�hX�6��u����*�����}Hg�͞�;�Xݬ��3!���p�Vrk6f5ӱ"�~dȄ����ۈ9OFMu_�Q���g��3s<op�d�T��0��/u8	����F6+E�m��ܲ�?dܪY36K��g���hz1����?��Βe�,��`G�w3!R���pԽ����r�Ĩt6�9�׏��p՝�`Ne1lĈ�X��~��Nf���n֗�:��b�I�?��8s,ֺ�ek(Ǎ�$��eG�9�V���l1��u��`)J�}p��V�c&I�(u���T����L�:0p���r�D��\��t�M���lF�۷�b"օ����qBj;P�PA��	�, h���0����Kt,@#i7-A3q�ВA���`��^�O٣�R��d~����vf�d��oYڇq4jB�Ί�9�l�$� �_����B� 7+H�)pJ��D	^�/*6d6�\���p��f�ϊ>`�ul~i-�8�0pV�̂�Q8l�t�g]h2+m&��b=�<ʲ��xd�p6�bbԤ2-\	�"�2n�fK`���Y��R����Uϴ4��6n�T�/Wx��L§�u�g1�v�V�Lү(uKS�i��Y:)�W���a�G50��̝GC�M�k�f��RD�&b]��&dؼ�lG�ם�n��/�jhV��8��b�Ь��[ⷺ��ЮǢ[G4rb Ḷ��~w]�������pb��,����)�_�[�Ac��r�$�[An܈Y�e�ҝ~Ŗ��#��n*��/疭9o�K��r�!#�z�K7b]��_�.�ɦ&<���h��Y�7V�O2�kON�n٫Y�k(f�e�u�r�)��9ZĲ����.�}3h�G�ss`7s�H�闘3��R��Bs3��Y�e`�L��u]38'�F���{�#n��܌��jl�|6Kb�V0�s�[��j�0�~�hN�u:7���U󆕌���x2.����Z�Q���>��s��e~��D�S�	��@	B�'L��,x˳0w��\�QΚ�QS��lz#���3f�)�Űy�uZvf*L���%�౹I�"����Z�l̰9Z�1��]��N��`,��yxp��G�ʩq3�����=1�[l5�8K�lN�D���!s���Ŧ"�3�8�$&�n�j��F�\72�x0dl��M1ud6uZ�s��k=N��j$�;����2�RNE�M���[�ItE���d�i�O��,V��U�#&F��|��O�sl�Y拋9l�u���n�@�FNĺ��a��wzʩ,��ލ�u��ѳ�i��Ì����H��u����#��l��3xYh�$e_������T8Z��� �9��$e����U�&1�^ٺUWs`��d��V�iu��1�G��s6��>*�as�Ίj��!�2�
���B5k0�b'b]F��y�y�:�	Sz4g��%#�����}7ɺcc5ΗusS�c#g]�,9'Ya��.��D�f]�gR�(uKe�.ڕ<�oC"��W�zV,7�o�f\?����޺��b��D���?���9l���G����u6n���8!�(O�d��� ��я�bn{zoFMi�sݸ9_Vi}�d�s��$�w5׿ʠ�\.h6�D��s��%�fI���Ss�.�c� �i9P�"rܴ򫰱����&�s��L����,7cw�n���yJ�U�17l���N�Qh�<��C�l���/���� 'I.3���r�p
�.�M��ڹI��МK�ڌ����]�e{e�g������C���$��^D�d	����ujF5lN>9͘�ds�r�ĥ_�����A�U%2+�����H���v���W��˳���$��
8�9T�)Y�ŷ�91I���C�������:�6�&	�;��9�E���ր����$�gđ6�i�����=���EK��
.n���z��$�~���>rF�S���ytݿ�W�A������ԀY&>�b|c��`�ﺅa(z^��6���j��O�f������9`^�$��^V� y��sbY�~o$�1+��r=eJ�3�0벒qej�	l��ӵ��a	�i�����tj�*�i��h�� x�� S����\'6r�j�p, ���w��䫹jn��n���?c|;�ઘ1S��N�2KeL�A6j�W�M��
^j+q�bX�$N�M�Y�5<�Y�M/�ut3 \�3PsDE+�&?����:TR��L+�i��w�^v�sG�G�{�)`��K�ul���]_5U8��2;�ǳD��u򮏜�����!j�M"bZtOr'M��C���I
��ɌZn��>0h�6۫�M����lj�A�<��ĥ�fN�C����c���Ks���lF3��p���^A�q�L�p��|�1��o���$11T^�W�]�R�������X1e+�f��2 P��\'0pⓇ��I:]�fΊ#��j�Rs�����sά��u�|���J����3��;�w�ʼpsdĘ�!�&Vi���l
VЬ@1h�l��qT^�{?O[6��-Eǅ���h�<�Mo-���-p�;Kwx�����v����u��ZĤ_٥�fY�!S�6��hο����鲦��F���:4h��K5N�5ZַMN�j`;K�MVe�������������X���Ǔ�0�}Z��r��!�Nҧ��J*H�<a�d���.+�B�����v]���q{e�,��f-' .�����B�Des�����RD�%&z�p��s�nu$��#f�
G�e�sb^ v�:1�N̡f����ul���QN����FO��!#��[P�u8����&�ʈuh�#n����������հI������)[�[x(<~R�x٦�Q��nZ�;P�Y��%1*�;��CM�f�M���ENL�M������u���[�ݍȉIʯ#����k݁uo@LR��Â�x����L׽�#fӧ`2������ԌN�pA[8��,���,�eh���:�Wj� Ŗ�؁�f���[�UX�#jm�$�{Y������΃���!ű������􆷨V������G�6�:4�se.������:��<^²��s����j���w����,5l��EhfV ��&)�A�f&1l���Է�iьe!R���p�-�Wm���$��@��r=�_��p�]ލ��:��.}���猛�0w��׉�`�\�lVd���:8n����1I�4�O:1��|>��4��J�:5�V�>��ob��90o���H��Y���J��~���Ix8M:����&��ު��XD�S�	��@	B�'L���"�0\.хf9,�Ÿ\�����4<��fj�~o�7��i��>󖑙�_��p킾 �7��R� -˅��߷$\E�3Z]�#�|6wwѻ�__7�b�#�p����)�$N���s"ufȜ�|o*���sxd�zlnx������]n����Cf!�ru吹��#ӕ5�jfj�%��Y���$���ʯ�!��*�9$��J���[�l_L����Eι�7�Hՠ��9&ࠩT<�p���l1oth�uP�^���F��5)x��}����{�������4z=�71ˉ=ulİ9�as��Ĩ�쮃0�s%�D�K9��`�x��y���؀Y|�pܴ���iwi�Ac&U�0F��e5��LŚ��z����:Y���8^��z����4���f���r��*w;p�WMҲ�����h֧&?M�ǥz�R~O��&s`�Ժ���<��I~�<��b�TN�y�۲�M&Fhfփ�����.��6X��D�)=8l��9��0[�7c�͏5BG�����r6
�܊AL��e��/�R�D�S`.fF�7�Ю��Z��}דs�#�b��`:ba"�z�-O4r܄)�*��y�WH-4��'�� G���f���cf�V^�A�0#1h��O68f�Y�j�S�@��
:�O�D�:b6�`�T5�QŰ9Lm��)��v�����&Y�� ���+f��-��|�JӢ^F�a��9O�,3����Yvf3x��}�C�b;7�k��،A��!#&Qw�Z@��v�q"u��l7s(:&��j6�c8��C?1Wc]�Y�ױY.r�ԍ���C3�Hc�HS�n��b̼Ne�2��J\t31�E�3cf���o����S3�X�h��[o2p�h�*5	����G��q��.Q1��hR�z�!����1�߅��03#B�0�ض��t��G�65���5W��h��9�ѥD�P�:6׏��<�5��3+p]�� a���Kv�-��T�_F17w����pM���ױ�f��k3ɺ��bn�6n�Ժm�fNf5p�s�2cf��x�lW�ΜQIn=�a�B�\[�f�+d���x'�*/�[������9���x��ѣ<��J&2#�
]~'q2��t�>�rYj��.�p?�?4�bFs���B�Z�m�6�:5� s��j�aS��9���[`�j�@7b����|H+�21e�/�,�b���u�İv_o5M�m:���3���E'A��I�~h*0�*�.lf�uG�ȼL�T׷<i��]I7I�'�a�4��*� '��s�I�,�C�5eS};P���jnb�G̒]��I��9�8�,T`��E�dJ���ˑ�ɷJ�Y����IY9efٯ��`��� (�
��$3p��Ϭ�Vύ���CE�5���p�N�-���//3f*��,_0�:mr�}�[V��!n�Aj�,_�K��]=5(�M0�y%�JxA=���]��S����A�$X~�����tUC��ThsܬӲ�:P�PA��	�, k��9�pYP΃�ԅv7��4`fΗ��L@8\����x����"�.��\�V� /p��an��$�r6W��cFNx�ذY>_0��D�S�Ĝ)h��ֱ떐���l�\\w5p���:����-(p���Adx�5�nˤ�����+����蚪9<�w��?t{���/��Q��V�M˼��,طl��y�J�w;��-���h��\��ˉI��;��5^B��8{&4��BL7'0d.�.\j`�z�q	�~�9��p�C��-��s�E��Ӻ�,y5�O�݃�y�]1j-|��C;8p�x5K&���m9;p�I۾�s��p�I��\^9K�ymx�t����
Oݹrnz�n���,d���d�˹2ME�Z�s>�YJ��u7�"7�Y��j�d�T#�]1p�3�@6Gw����5��T��H�I���9ƭxz4ci�ƪ*&u����c]帉�����z?�9a+�4[�u#&ja��|81�98�K������&��͊���R�Ŕ�YS7b��nn]�MN����Ϋ�ԉ�v��.�ڹqs�7�$u���,���,i���ΓBN%�B{0?Z����n��b\�[��b"օ�'��qBj;P�PA��	�, h���0L1'�%:���Ҵ����9��7SC�����E�mR�n�_�$�^���ަ&4��䐹��%	�Q��VŘ�=�^ņ��U��M��'�b�#�p���˩�$N���"uG[��@N~�&����cs��U�̦��r[�5=�51����!#���g]/ϲ���\4���$R��Y��l�d�U��Y�Ko�W�L\��es՘Y��u�?0��Ax���&鯞4/:��N��U_bG3�/`R��X��bހ���uL6Z���F��e5)��l_��q@�d_�u]���DL�ꂮF�z�Yn��M[w�d���YQ91�-��"��\I2�RΝ�b/�E�tÓ~�cf��.�v3+��{g�&u�J��͆�b�u+t[���S�_����r���[�x��OOfio|ag#��V���%s�WMҲ�g���mM��K��ȹi)��ny�ֱ�q6�n�9�nd���&i�!t�n|[1j*���s�oxi�����`���d�E�����V7w1L���aCF�9�f�U���!x!��W|�¿�Kk�+B�M��ԭ��o�4�/��'����d*�̬!5G�A<�p5�"��`8Z]�xn-�������%Z�Z���N38r��)�6��+ffqW���*����A�L����v2�l�}��!G"9������.2U54�6b�F6P�qBj;P�PA��	�, �<� ���+f����j��%����b!��@�T�=�nb�[��4�̨�^bpP%��=�*o�V����p����#�����k���ɼBn��g0b����Z/k6���R>�9gb�f�WyI���/0n"��n4�Ub��@͆Mxү�mZ�+u��T׏�-ќ�j�Tg��
c�_���w�W̉�LG�Q�6j�\��*0�w2�p#5�&���¦R�] ��[.)�&�R\7�����n���I��f��l��R k�cfY���Xx0^O5K�K�+8�W�r�,C{�ve=�#�,�Gm����#1o3�d�ԏR���-��smհI��&��]b��Cʺf���n�\Pj��[�T]�kz]��27p�t�>"#ց�p|�ʹW�Mx��Y�|ߺ��Khh���ݯ��,�Um���9��I�f7�p�����n�!�f1nǃ�ګ��{�g��� �`f���By���Ҿ�I���zƃ�e��QO&L.�1<u�.�I�b	Ɉ	S���u!��[]_A�����S���d�i0IE���b��ɐL��,;���@�����첂C����,�j^�,�u�llӻ�#,�Wf���#�j��v]A��r�Vb̨A�6�ͬ�!�ps��&ght1,9�nח����Y�d��!s�U�.�_�w��W+���D��w����n���Huh�l��ͬ�����Q
���ġKM�N��}��]�&����2B#'�cl#k���� �.��s��� 4�I��Y�0E��-3r��Qs�-**��v�����&Y@�s�}���(��j��b�<�5�IΡu�0s����0S�oz����c���f)�	�ug͡;�}��tr�VN���,8j�;�d�u[����z�-ۍ���zau�{���
M�7�,�ܶ�X�*䘁s�9��·� �YWq_L��pϛ%��ĸI�'�@�pz��pv��!�L�"՝h��>�$��Rgfp��j�_�d��o��#��jݎ��uȌ���|��Y;5p"�e�Nw9���r��'���!F����Kq��9/|'�.0����`��n��9�d�İ|��C.W6�x6k��o�!N��tY�d�lzy�)֭ҢG�h�$�O�%Gf,����X̙�İ�uS���Y�ȃ`޳C�Ll�$�X��^�G�a,b]���'g���T<DO�ู�nf#�:� ���A�^�}3����J�`��yx;ݓB�T6�cny'\�T�l6�4t���_��)�B<��T��-q31l`����V�s�I͈Y5I���bZ��ذ��c�f����0n���!y��1t���������J���'��5g�fe�3j��)��v�����&Y�_�z�Ჰ���vJ��Z�a3�4M�Z������~@bf���^K�Z�+����:n�fy���F��hu����\[8�$�~�8�o�?D��7w[�f�$��c�
gl�3\݉�fo���c3Y&r���^�LksP��s�<�׹z��:8`�z�{��/J��-�$��n�u��sd��]��鹿��ڤo�c�46�����<s����ub�G6���q��Q�&|`���뚀)�����O�� >��w����r[釄�T��eC�R#'4ʢS8�}��('�R3���qs���f��Z���p)r��h��%͋2�NLX�Ȱٌ�E�,�[��]t�E�/̂#&(��+�͸�#'<�_�uX��6�A1�R��e�5N�N��%x��d�Y�g���I�23K��j�y��l��Q3�Qjb�n��򆳼���X��[?9(F��%)&<�w�,�=6� ��~���0�iQ�R���,��!���$��R��2�[��d.>�����6aͥIv��%�f�Y7G���u�rC�f�ֹY5��oɲ�f����V��RV��ˊ���,�f��lȼv���b\�dF����@� 5`V֌��Ɩ�" "̐`�LB���G�a0w��6�Vjج�f��I������jĄ�����F�72M�-%8`���l��qGݝ[��T���X��k�Ÿ9-���$��n��A�ep�|Z+�2g��5�&b]IOfY<�ܞ1L�oӱ�XW�֑�RwW9I<��L6�jUИ�֭��n��5K&?��U]m7շ�Y�<h�s�e�\��pJ���9\$��+���S�/t+��_���X�f�]�hVMu2�s�l�g#��ݼW�����RV��b.��.<����4�2˙ ǃ��c�V��ȁ��p
����l��Q9J�������7�t=B�*�Yb7���3�o3��us'̸麕8��L�qR��h���ÉZ����P���,�%I&L���z��ԡ��3����d]0���I�f�a�;�
d�j�º%ܿ�r�l�M���<$��q�]5���h��,����Y6b��ݰ/GI�b�&b��nbd^N�� ���.2�����pxү��C�Iuȭ|vs��̜N1�7��K|]�/�/ �qޚi�̩���Ɩ�B]E���� T�~y�$ȑ!�0\��}j�b6��
e3Q�iSG�ѵ�Ade����W���ܻ�3՝̀9ਁ�F��$?���b=��~1f��#=�$7����֧�;6.��c �[��r�V��oI,��X�C}R�u����q]���d�lz�Ȉ�����H��<rِ)�[@�d��M���Q�{���b����7��O�#ee�/�9�$<�n�	X�V��v�W'Yw��iD�j8`�_M�70��]�}4���j�5WsBI�fx����)�~�J��똄�Hu��̏��/�nq�z7�J�I�+R�z��+_�&���T;|�Y���̑���^���C�6���攙�|�[��N��\n2l̬;�*�0ԝc�s]V����
ss_|/I����y���]�|��ͅ�vquh@��ʹ�d���ظ����_������R�0�͠:I�3�8(����w��fuN���,���udƔ%��N��m�������X��7�U������N[6�M������\
r����`}����$�#�-$l䰁�-r��^��fy,�j���Q����&I�3���:7f*_��������}8��cUN��o���@URhg�1g��u�z�sڙq���sIͭ8їR��ͯ�w��P{!]G1ϻ(��:0�[�p��e��u�/9����gf!\��#6fj�W�]��$�O29���ifU�D�K�L��!f%�Tt�!�BB�a�e\ܿ䛸�K)F~5U�k!DSһ9���,���zV4/Y9r��68n�^WM��չ�K�Z��}��j׺�̡f�Ĺ��r��]4��g�z�㵋ᘚ��n�e6�n�~�K�]hb�^���=犘j�
_hV�i�&.y�:6`��V8�^��/T`��[t�c�G�l��1���������L`��d"�e����.���0�_V��:�æBӱr>�؄AuXp�Uw���\@f��qBj;P�PA��	�, h��~��������"F�T!S�6�H�_��n٘��n���qx{ŀY?1���j�]��ݬ���`��9�X~lȜHhb��x���s�i��Y�e�Y1)N_74Y׵}��2��M��H�~�!c1n��QNĺ���o	^4+V-��~�w��mAs�����0>��R'�@+΁Í5n��E�[�`��S9��+�Z���_�7��������u{*55�e;��l�d��|W�]FH�]�Z�Y��q��G�����w��Y�k��ȉ���l��ȩp��G�,%6nR$��]���mf*����^�hbe�R���b�DN�D��.���#�Ŋ�jcn��;N�l��9�n�ě��l@[�J�sh��k��^ͅ �6ɺ����!�.�y0t[.9�I&o���_pմe�6�u)A�sᬽ�44=��W��]s7ɺ5;�֓͊V-tl�,k5r6��%9dO�M��j�p��7r�z��*���9�Ԭ}R~9k��0�»p�dS�E�u���V���.����������r���z1ſ_��/��SMQ��O�3C&ƿ(uKw���1�;P-�_j�� h��,�C��$�n��a/8���uYx`��3�����bN���+;��P���9\H��-$bNw2���B��cN��u_�'�3P�jeօ���`�_�g\5n"֥��sO��=<��,������]���Qg�V��(e��M�-ih��e�8�l�XHb8�f�|ï��M�B���n��ac��v�Π�u��ֹ}��aJ��d��Ä���5?���&�K3�N'D��%�_�0�r֊�̊޺E�F�Y��djӦ��2\�m�,��_�|��a��sc�Ll��|Jrs��|pN11lB����]�K�ɺ#�n|Y��Fmd3h̐9��$�^���x����E#�̹}T%Ai����oFMĺ�߈{8!s��	S����ȩ\���R[]5I*-v7d��g����B��y�`]�����Y��޵J����Z�~��Ed������f����~�Wc�P�nr�	Sz2�|h^�j�}�n(��'7a�;iΉ��"�_����ވ�3K���-�m�Q�lh6f���7I�eK ����@��$��u���Eu�W��Y׳Nκ����y�`�q��,�����7�P�ȼz��d��2r�.�Ӫ�Y&d�؄'�y���Xp�7��;�$����[��{Q�YI8I�D��.,6�Q�ƍ0r��	��e���̦���L�S^����y/��*�pf�D5w<��͜Mn���_Y�&g5C751���G�=1a��g�,Ni2h"�5�w ��%MT���p���'?f�l�qѠ�.<ed�}S75�ND�����������
�+��v�����&Y@�,o1}����y����2�3 P�65@�f�G���035�
SC�0���d��dj��5��s����C�N�Y�f�/��.&Y��E��%x>V�6�����$�_FfKp�`�T/�`�̺.75I.���񉸌�D�+�m�	�ͺm(<�w�20/Ы�ùx��&�y`i
��Mf�c��#��ai��T��w���h��;o12l���g�����_�0}f�q��6[�	Oz2p�e��N�B/5C�M.f��:9�'���q��/J]t�.���� "u��͉6�^�IBG�;�,�n�0bb8�����3p?up�����nhĨI�G��R�������ʘiF�1����CƲ\f"���j�ĕ\&+M&L�ټ��^DO���Z�֙ͭK�?J�ͭ��3��J!x|]t�]g6��j�YJa���e���Oa�[�� �P)�����/$�Dہɜc�f�]��DLr8'���V�r��և����d��6��'L[��e���j�	�od�u����Z�ӟ�ǃ6+�&s��b��ф��̺������$��ԅ��rԐY"˅1�lE���� T�~y�$��]L`���p�q���,8���(8���T+��/ fj��,�3�� ����!@̀�&��rK����0�]�Sr0�!��z��$���Y�Wm{�Ą'�-�-l�l �4a�[����]/h�0���r���I��j��n��	ߖ���1���3a��(�?����ɺ���hV�Z�ɿ��b~�y{2a�[�W�|�	��&&�Ɔ��%��p��[|E3:����Z������xv�@&ȊZw���ݖs`I�w܀Y��6�J�9��58�)e�\S6f������zɂ0�Y1uh�,ϕw�Q3590����B��+B�9�f#ǈ3)c_&�P9�B�Y0w�
-D�2���d��L3t�[���<�$�!8f�|�������P6��/���!xԺ�,qcf��Y��:,P�.:Cݬ�zp�Kab��m��eB����X7p������)'<�T��kB�@�L庪	������GMu?:��³<N��uC&�1|�޷`>�Nͦ��Y����	� f���q3rB�nsf.���$�#�]��Z�d�$4gfs�u=��k��](ce��ޟF�7c�����w�M�p=��w�x���d�qwd��Fj��R/�m���6�_�S��)<u��s�I���y��<<p��HuQmL2�r�-��JB7���|���ń	h�}��if�(�Jf8��)��	���*ll)�HM��BsxV��39Y�$�s���S@�	sUo@�5g��'Y[0+�EX^��@O�~���G��,s/�hkj�LҿHu�:�[��;�_�:1O�^'������oL�8d�v��/2�!u��� �%�dl"�e�-�o���j�͡�̊ޕ��ٶ�&����ues�VM���	�[���&�է����uS]73���ͣ�������j����υ�?��ݷuz(9��t[����{#���b���ֽ��Yć�a�=��ی�g\�=3b"�eN���a�pO&L����J/�'�~�[��g�n"�u\���ub�����|�T��K��r��J����or%F�IՖ���pF����:9��J��L&���_2�+�B�aqo'��U9�VMa3��h�3,Fx'��Y���u��e�fyX��uE7�JfЈ9�u�z>��:��������r�!�L'D��%�_�0��d�W`��9����b�����uӦVsI/�mŜ�fֲ�>�Fw9/,z&5I$�9Zݬ٨+�L�V��=�^0�$�6r��.9�C��/��#�0���tY�$�[��d#�$� �u+�ʠ9��I
�P������
�h���E���ԓu+�±�6b�|ĺl�
|�ö����d��]��� Y�����lX��$�G�;�ݰY���+��E�CsX�b����p�&�%#G�`[���Rk����̳�Gr:���5�T�q�&N��q)?��5b]ʱ�������fѬ��7��p�ֵO��Y�j��
5`���A9l�(2I���9�$�t�2X���~S���!�S�f�����x,a���S��T`]�rkGN�>g�4�v՘ɠ�����M��G2�#���iҐY��5��:6�&����z�!b]��D`[�k��b�С�"���9��!s���1��Rg�\��⌏R�����ߓ����ݑ%U g�3�}���9z6��n
�Ɨ����-���f�V,L�O%4&�,G��sډ�0m$Z���S���L�C�F`�\��&��� �+�rj=������z޷�fUN��f}Y9�7E���� T�~y�$�AUL`���s��`��y���f�rNh�ec�_�`sG2�CJ���Z�Ac<7�N��i"�L��-��~�M��ki=�Rf3X���q�lKC�a8I��?�&��U}#�f�fdj�$��\�U^�̀����N�wn�3aJ?(Y2�rj�e����:��aͺᬒ��̈́�h0���M�i ���b�$S?���"7p��	��+�)���M8V�e��Y�����\?2�H��͈9��6EHj�rw�i����\���$�0Z�����g��Z����9��	��e��ͱ®�$a��F�lr�X��p
��r���Je8�zn��&��V�`6�m���:7kq��A&������6�.�_57��hN�0�7�[x������ܺ����ڼ�X�nz���� <8j�c��I�&D�V��
��T'�i7o�������AL�&�g��dαA���a��İ|�:�^��{�s���C_5��+�T0c�He�&<B[����
G��m���<��u9�琺��2��t���SFfݯ/0jԠQ��T������!����Z��S�8!�(A� ��I�R�`��B��̜���iS�jVn���|����p��Y�_6���k�x�_�Ź��`3ٵ(un��;�v9o���V�	��eG���]9�L���.�i}x:ﻎ��ܺ�	N���6�F[�u]�]g]N�5}KL�f!��꒩u�aͅ��!&�_�����hШ9��$����,N9]w�`V�'�[J���n��r�]�G�/%��M��A�������lB����D]K}�)�Հ1���z,�ųd�`��8�p�6���<$�T��%jm������N�(vF����T����f�._2�U����x��,j�] g�,#2b�晗4/J��:1a�[Nrڋ��d��_���!�x��.�uE�lpԀy8�}}ό�oPL���Y���Qs}�r0K�-�(1�/47}�48k.'����`ج�";XW������ƨ����e��e"Mĺ��z.�=6�TMx�/�eww��ZM��Ԉ�YG�p�mnU����M����p0��Vs����lu��2d�`��Huʹ��t7I�.40����]�&穹�gNL�B�f��@d��엚es:������K�_�YG9�e9��y^8a�;
W�b^�mcHWH�ED�!�����+�0�a��ն��3�X��5p�0�F��bl����G09�e1��Q�k�.l6I��mٰ�f�l�!㈸gw�L�\/Q#��J-�`*C���Z�����9��m��!�&b]I�{*^��Ô~cj���@)[�r������uEg�9�T�.!7fԜ1�ϰ�o��S�o�3�͠i�ϩ��pSRo�B����dݣ����M�Sy�/����b�+o�����6�F�MS�&Ff2��h����KY<���!INx��As�ݱ�FN�[��n�L9��ulVՌ�n�BS�sp�W�Lu�ԽL�hpJ�I��βXvj"6��$��
�k��K�-�l�u?��ᔜ��v����.���΢۸7b~Y�q�f�/~8�N��Ŵ���L�.
��>n����ha�[�dN��yF�Y�����6����~�z�j�ġ� a���v�BA3�g��I�g!8��_N׹�P��� �&�D�v@cfY��X����Ey4�Sx�?�R9/���z���7���`k�u	�1c�֭˚t�4���bn͂z���Q�	��@	B�'L��9b� sT���f�^�l&�4�dwe5�=Ȭ35���ѹ�����LugM�l#_@�$��t��ǔZ'f<Ҧ�/����
�9l>Q���.g�O�$A�����j�1S	�4������d��?��.��>=O�$�,�տ��[�b
RWY�%^�bӯ�������N�s��ރ��pA�m�舶���	O�;���fdȠ1S���r�����А�[����{��uj����,8	�V�zb�ym-��������2/7����н��똄�(u붜wɜ�^�o�527��W��_���H=Nυ$�Ŝ�hvH��[��#�\�1e�� f�k6fȬ��%�2�
0`FXa�[>V0���eR}[�ͭ��[4I��{p^��j�����غ5]&�|ܡ�e��T5���odVv���SS������KGX3Õչ�5�}Y��Ml��'
0h.4dj����Khy-�I:���-9�D���W�*.��М��I��Eq�9�n���v�Y�')�0��\��+f&��Hu��f��r�T&sXK�8��uw�h���l��]׍��j������ts�.�G�a-1����5�՜�1��)�zp�g9C5as$$�eӋP�e]V�hQs�Ш9^�Qu��2=|׺�ssN����N|݁p�%�6q�����j���񮮻3I~�T��6l��5��"��^fF�4aJ�2Ά���;S��g^Bl�S9�rZv�"CS��9{Ԝ�h��ʅE���Э�
�#g��@Ӳ���Y.l��&������.����!�Z��ׄLK����Ĩ*�N2뽮ۀ���i�l�� V��=��%41г��,'�����,.2�p�Z���6{��k'�ߑ��Cs���1����$3`g�b���:�˝͑�.�w/׳�u���p�<��r��� ��3!l���j��ᄫ��1�2b.]�"N�@mJ*H�<a��V�0��a��
?1��t��9���v{����nN�3{-��0�*8^v�i3�GN��uK�ؖ��a��-�l��ZM\����"X=1-����˱���a�{ҁ���FM���c��k@f���`)��d�D�+\_9��:-�p�e#�����d�Of2ϻ�$���sTV��j������c�/��o������ܣ���Ǡk�/�E8H����
K����������i��<��ڬ�6ɲ�.��}�����2��U�3tZy7�I}�J�ɲe���7YW�M�Ԉuh.��]��N·(u7����h%c0�t�"��u���-ֽ��CM��͂fA�3�r�u��;��Ic���ԗ��߈u)�ň!��s�L8ҿ�`~��%8�n�Κ�;���\��N���f��zg��afQ�q��Uq�����I���-�hVf��
$�_xlF3f�4ظasl�Dh�N��+�fQ]���Z�9v��iyÕ\�b>f*���IvX<f�I��D�Fќ���+l�nVb��#f��#��pW�*��рM�����؜�`&�B����Eaf0����]X^�58��Ī�v��x}"�e����,��*\��I��R�S!��2sy/�s���dws:\̈́��ƃ�:;͠���%��|g#��*�bs�`�1u���wK0b�D�����zI�t�#}D�/�So�,���)��v�����&Y@�H3r}�B<�e���Ԧ�x]��yї������1�b���:\�vm�����亦@��n^p�Vz]��	���4K�!GL���Θ��Z/2WW6`��Z��W��fk6�n=�yq���I�-�e�8+�F��uٷ��6��=Sz1���#w��aS݇soĠ9�����g�V~CnȰ	��l�r�V�+:,g7���<O��2�U��"p���z^�������"\З��l�'����jb�Tˎx2n6���.,e�z�fsR/r�$��+�<�e��r�̹l}�83���!p�ܜif���7I�Hu`N�[�	0b� ����UY;3l
Ȭ��k`�&&�Ȁy���9�Vز��fbd���0�r0l"֥tB��`g,5�I��?�*�%)�M��ln]�ߑ���:m�f%�$[�LܐA�x�"�0�?�n�;Ȭ�c|�:0w���Ԡa����/�Q���ԡ��2�&��u5���4.������j�[�j����b6~VE�wZ���D�&2��o��ew[�1��	8`�l|Y�ɜ�͉�0�	S9h��M�YTnb��-�/�:�Q��{�.E���� T�~y�$�B��� ��`��A��´�R6r�ԦM����d�KK��Z��j����.����r����*��1��f��s�	���`�1f+1ɺ��9���E���YBd6���Y2IF���Y�p�o���X�j��V���r5���XV�:���&ԸY�e��g�}X"��h�I���Z��^�E�Q8kG&<��q`#�FXΧɹx^$�ߊ; gӫ�&L��J.8d̬�0�pF-�7/l`Ȅ'�pb�n��U���͹��Z,���]���HK}�n��ׅ��^}1n�.�����[�9�O�ő$x�:0j�[�90b����0h�P���R@κlN��nL��dz4��M�a����:8w�8����_͠{ebd�D����8u1aJ��u�vb�)�;�n���%��n���:m��I��ՅCx�v��p�������< �	7b���̝�cf�M�I�ݗ�
^pݸyg�Cg`���d�!x�����ȁS9��
^��=L2��Ӹ9}��15��,����0qlݗ�:ޗ���u9���҇������8B�0�	S����`�lha��/�0,|���67|�p@�"N�@mJ*H�<a���/�0k{о`Wsu��r\%2�iS���+�=��35��6g��9T�aӚ/�M��^�$��j,��.�+�&Ludv��y{��e�,��l��D�=6�fA��j܄'����]���b&Lup�lJ��j+�7l�\țT���	r�����ï�~U�]�&�b��_�����M�ͳ�ag��Ô~�ٸ�6b�0��6��k��M�D%1!G��F�f������r�r�������Z��趿n��9����br�՝��o�ޜ0�����\�[_9]wM�kas3ҥ��8W���o��c�P5����24�x-�3%�z�Yh�5_=1Iߢԭ7�U����Iԑ��|VeQ��0��Z��M����~HZ��Yh:�bZ ���Css�$��1���9�����n�N̺�p1a�.���`�9�B��@m���~ۺa^h�T���跹����/f����is�fu�\��?�X����6��,�s�������uցQSݏ�p8����[ߊ����u��f٣9��tp9��f���QM�o�}�V��{pB��_�l�%���$�#�-ݭĜU�]NB��<��1��C5�����V��X	&�p7��+�0����s��9ߖa��uxݲ����H֑!���^�� �����(�g=��[�'���������s2�I�e�0,�%��Mx�,���0��d��ny�9Q�����f��
,�j��	�F+��ᠹ:M59��P�np�$��}Y�Y�`�1���C�3{waE�$떣7��]�����dnL�ej6��.���������y�5N�ߌ��F�´�6u��x3�'��T��,�g�&��Q��/J�*/��:��4���w�nsɴ�pĀY��,���-7~�2j"�e!n�_H[\���?�*d��禸���v41u�uf����l!���1�m�� {u��\��C�: �����T�V�����&�6hРQcF��Ŧ����,�`�\���;(ۋi���Z*h&b��K��*շe�c����`׍�0%Gs��W�Ku}ŏ�M�a3&
����F��t�?�
Zda�����8��Lҁ(uw�%�Pc�[^��/�}�o���*�Y!d���ۻ��ח�
`�,��:b�Ġ�!�h�>�8h�c`A�Brŏ�1��
f�ͮ3lb���4���V@\���t�o�߲\x�o'���u�8!�(A� ��I�%�<� ���}�s��Z��ڴ��<��ː�J�e����r_RfN�J�S*�D3���0b�]p��=YW2`�D]o1�8h�,8�[�����%�s{w$�C3	�|23�f�)��瀙UR��z-9ی3��l�������;@��Uc�./G�}Zo4L�w����3P�urH�as ��-�f&�I�ʤQ�NГ
�B��p���\�]����]���P��I��z�9���D[�.3�%1nN൏���;��9ƣ֥�Z4̍�j~Y�9��,��#s���f��d��e�����V�!��l�aS��R̘�:�iuܰYo6�"fS�|�,/6��@с�u�%�8�nn��v�� �A��}N���V�(1�V���1F��Ux�%ܤ�st�Y'5�ঁ9ֲ[����h�D��������͘Q����p!+i�"f������T�n+��8<��n=���=n�22p��ج�����Ay��n�ȉX��FW�4�2L��<�ɸΗ��?�� ��01�������t�j�_��7�LF���-�al���ˏf���b�8��i�_��Syp���Ż��V�	��@	B�'L������([�j܌��`�?[m��U%s��_��Z���U9��:n��oԨ9��$x��C�W��*u���D��M�-A0d�\�aaס9�։���|�p�+1��ӧ���vcf#7JM���z<�-�d������esF/w7d9w��oU-�3n��u]�q�f�,H���!LƋy81+�up��,7'q#*�~%�܁����&L�Y��z'���G��ut�Yfn�������:���dS���P\�M�n�ԭ��.�;�@_�f��,�s���Y=0lV�0r��څD���03�_I�G�[j`��J3��$������B5\�zD��ɖL�Y4Ǜ��M������m&��G?��\`�D���R5��y�,'?��As�Y��da-2'V{���^����C踺�k �`sD.�����w2�����̝X �Ss�Ā�,�Mo�uh_�ҍİx_�|��a�N唛�Ь�햩�d�U߀5p��S�Gh�s��1�nr
G�ԥ=��Y���L�8�*�>�ݜ\)/��&Led�9���Y��b����-�r̸!��̈	�qBj;P�PA��	�������ڂsϗ+�ڋnYզM-�stEo� f&8��g��[^h Z�p9Ζ��]㍙ɮE��~��M�W=6���EPu���(иy��E&��e�� 3��N]��#s+�W�r�ukz2�M���L׭�ZVOh91un.0��'#S��s����]��$��Rgf1l��1���uknf����#s;��u���-���Hp�T�OG3��{r�I�?ucuЬ�nt�Ga8�d�
Y ��A��zq%@k=��Y�k�FKM�ί�h3yߓ����[����(9���0��pBP��K��I�������4Cf��XZ'h�N��"�HМ�I������k�F����d��_���"�x�/ȵ	E��lpԀy8�`}ό��ݠ�)[��G�������ܬ�b�T�������^s9D^w` �f�/��N׭�f�7FML��Y�\&V#�e��sY��j|9l���]��|	�[�:҇�N�0n��Af- �-�.,�>�՜3�o�����I��(h�5u�:0�f�!n�V^�`N�忾`�n9�Y�S���jb�j7���G#�he�/5��tq���"<��4��Y�YG9U�u]��x]7'Lu�0.<jn�11���$�"(��d�LB��X�аy�v�_�&�@�5p�0�F���l����
G�<��v+^��-\��MR�u[6l�(���4d�����d��k�O�c�2Xΐ���\�$����_�4�J��Smy��S�E�f�޺Բ����&�"�x�9N�Ժ�ߍ�PN���$sF�j�D6`��4��ԋ���ݔ�+����dݣ�����+u�ׄ�K��L�U*1���3�A���n�61��iPXg39F|a��qb�mQ#�As�1�FN)�U���<#��lV���t9+��YG7뺽�8
D�[_8bF�c�Lҁu[�̮��9ɓ��f���;��t�ٻF�~�V�Q9Ͻ�[�0E�˼�mO���,&L�7�fK}��)uǷ�%p�,�db
��!�3�uZ�ٸ1��ͬ��.����%XW5��o��g͏��D��8T���⛫�'���2`#&��ဲ�wKN�]��.dk|�őp��%�,�D�Ko��J��#BMx�?�R9�,�ru� z�>��Ĥ�O�v#̘��I檭�����X�-Y���FWE'D��%�_�0�r$��� s�>��y�����t��9`����pe����7����M,14��<0��l|�V����q��VUC�l�6�~fb�\�����2�⺁s;�6���0��)����j�i*����9d$E%�:�S����F�\�#	KH�:��v�JLE�U73��&6���ݗv��A�X��q��r�d�57#��&#'<���²�pI���9����Гu_����֩as���5Xp�������� ���ڼNL�˼�ݬ�2/��3\�1	�Q�.��;�/��"�R��_�$�׉��`/n$�-�4D��Pj̘��W�6���&��a��n0kQ�.�5Z��N�r���o����l��˷�k��q�/�E����}1_~,dG��j7�����2_��M�i� ԰q#&�'��ؕsV�S|�<�!��d��c���6����m�Mof���%w!/�� ���,�'I�#�`v��ͨ�Z�cmۊ,��'L1��Er�?��)1���cb���p�QxJ�Y��l���Wh�����9u��=r�$��$4ƪ��:4w�کyW�B9K�nb�nr�7`VN�P���:��M�- d�p5gJG7sr���Y�|s�Y&as�&����˼���'�ew�8ZF1Y����pY!ne�ܜ���%�_w4ߖ�-\����f�g\�uO9���3I~�L��6l�쩉X� %�E�23jܠ	S��Y$Kh�d�'4w�Ms*�_N��?X��G�F��Shb¢���%+X��e���n.'8��h����!������.oH���M%��;�؈�a��yP�ft�e�x����p�[6�` �ҍ��g=�b�k�wf=$8b�T��4�p�]��ꆀ�j���aJg��Xg7fb��:9/����:�c�dY�l��hu�G3g����.pܸ	S�u8��9P���=Hql�|�Y�}8h�Tw��1�2+r�V�qBj;P�PA��	��5�`��9�8+fV�q2x��^�)�������ws�М�����[67���t�v��Q��<Γ��̒����\8w���(<�Un^�\ŀI�|ݺ, l���Twspo��&��j�\ +}����~R�����S�� �S���\����&�nqoZ�)}:%�X��1{�<���5Z��?u��[�\�7-���5[�5�E3(H�ml�뼚M4�y��k��_���yT����J]�M��������|����N]�Ɇ�ۦ��A�<��t�I��EO�Hw��;�/R7(4b*�/��:���!n~�'����J��V����|ݐI�'�fC�j��T����p�bn�A�Q��	"f���!�_�:3d���yG
��}1p�Ҍ��;��!�zb.EL݉���U�4f"�e�����]dj�zaH��29K�,6l����Ey�Ȥ�:6j.�&��)�����O�����s�nda��~�y�\���#}���[T� 196�L�O�Q� 	��w��{��� 6�``�h�#�Y*����.2��RΉi�$2r|�iN.DkO����,�`䰉!�7��iY��j�&spS����K̯������^�fR��ds�z�#�B��-�C��3/Fv1�0����B�5`�u_8�w�O*1h�7f�^�l6���hb�zhN]5�ܛ^rn��q�)���\��w-*`-g0K�_��o�\�ۜ>d�D�S�	��@	B�'L����b� �e!��Ve��Y,�i�[�6�����]A��Z��l"8�0�6Mbn�z1H�������)��K�����I�2�԰���)�s�����&I���;�l�h�SA�P{^� 5I������웑���w7��F3ל�0�?�wgǢ� �����^M��s�.l�u%L����]�2�V��x^$#\�����l&L�Y�G��#��u�?4�n���׌��_��7d�M忛�z`b��NΥ;Gn�J�I�['�x�q�lm�̒Tq#j�d�a3�����L�����qL�RF�R_��b8+���_8���Z�^g���!&	��Pf�Y��hUT7��?�Mrt�b.��.pb"����j��I7aJ��\��c�æs�d�z-�$/"�������������Q1���}�x[8�`���9Ԛ	[�q́YJh���b���r:�2'��Ԭ�nL�ͮ�C���M-[��KF��M"9�����5Ta��p.ρ�MT�R6�n]/8QY��_��aŖ<����4s���v�23�����:ɹ�����R�Cκ�Y߰@�"N�@mJ*H�<a�d��L/��ո9ƥg�䐩M�#���+w�]�(f���u_���_�����&���g��/�nf�Rw/�<�
'~�}U��+�nkMF�FMBf�O�-�����Z�Y�7LM��&G�`�}/b]��:,39b̬dE[ғ����꾙�x��k�����T����R��K�Zwlʹϛ:o��9����߀6�q�̻��V7j�c<��S7{瞙0���Qs��(�����o�ͬ7�;�9Gn�J�I�[D,`�,�#ny�	����e���{�K�B0r�,7d$g�}�����L�[��|�ݘ��d��v�����f]��H"�@��_�h�D�K�jf�?�זLxү���ܮ;���Q2g�K�$Rݡ��&f�!�_l]X�y��j��;�Q8<9P�|
[�r(#G61��f}_�XVSL�(4n�pE��D��w/�Ħp��BCF��ML���,�KR�0	��_91r6� St��!�̈�&*r��ܒ���xLa��f��Ÿ����r�ͩA�&�s�ua���[7n��Y��i
qBj;P�PA��	�, �1}��¶FnİY��-�ڴ����O�r$35������;�ڣsXl4�u0�o��L!6a�ccͮ�/n����S�I��_�`Ĭ����l�,���r��)`ݿ��Y?6p�T\ob�=:��FMLz6n6�d��j���ӟ�`�6�t�
#��By '�nT���(�}�0E���j/�U	���b�U'���&�>��*&�ʆ��e��k3F�i����έ�9!���0ؿp̬�KV��ၣ(���A�<]�lΨd��.�-�(����-�^M
�/ss���`���6�����<A�n�ˋ�A��j�z.�k�@nt�'}�R�0l���1�D/�5>K�e�^rɠ9ǗՊ�ڤ뷠�Y�p�~-��\4�c�_���m8�\�y��[�7h&<�����彌�{p܄Fa8��-ӛs�����a�Y=9������,<d�6�at���vs���}���`6���]�lVENx��͠g_+2A���ВYo0��L���ܩM���	�6�3pW�琨Ɗ�j=W��x=�U�F̢s�,2I��gd֏��Kp�u!9p��ʷ����%ј�[�.��3/gC�`��5V���|��!౑,\tKv��25�S��,�c0��uX��]57{%�2sŜkS��e��f��	.�9�0
�̀	A���7p�. Us��쯾�[������>����pp��*,Q2G�b[��4L_71k��ɜ�n�u�Dٸy����e�f(I�$Yyr?�����48/�њl��D�5[
�ic+�����Bw�b�a�[*��c�rI�������p����4�M[w��72���1u�7��^Dk�.��f�g�a�L����вZw6r�����V��:8jN 7p�-���V�_�6B�M��]��f�Tնg�r�	4qt:1��p]���A2G�D���S/����m��f��Y�`�]H�$�، ��Ȳ�ul��'Ǌ�����;��:ɉ\�r���ۭ���7s��ff9b�������ĐlY^2p�����R���0�ݟK�4��J����s�^�I���m�̒ �M��`edb�? �Y8���nr�̼�n�;�+�9G�����cs=^�&�7��e#ͻ�nrnɲRs�+�@�8�`�ҲYal�:�������f���^��"Pہ�
�/O�dy1}��̅���� �F�ڴ��\�%�����
3SB�	b48K�f-GId�Y0�x�mo&�pȸQ��7��!����
C�Fw�
զ�h�d���]3bb����{�d*Ա9p��h�\x�EC��Y������ j��S�<�f��p�u�?4�g8`VVM�ҏ0������8�[*�#'	���̬7�{���2F���ccQ�YI8�����1�0��nݷ��u]�a�b$�֍̅�\ͼ�֝"�k��l�&�����F�n���4�1�ba��,�۟�r��:2_�0h�u��̌�b䈩�kp4.Z4��d�5���P̦9���Y1�:5�y/�;Q�X/[|+�L\6s�f7H�G�s���I�s�o�x�x��nN.7+���8	VO�0�_M�0�����1�&N�Y�cc&b]��������f��&� �b�NF�eFs��TwT��w^L����j��y=lLB�&<���`�d��vm"p����.ja�q�/���7?L1�
�����R���d�t��Y㡹8�[�<��`_M	�}a8�l�rUw�\�ׇL�3k������lJ���ON�O'D��%�_�0�r���1([~'�`{�,�V�6u>��r�]8ֲ?��͢9�:8���2 3hN��M����C��^,���
9I���l؜ߍ��%3��s�Hr@��Y�W�gsh���/Y��.�Ë#&b]���/7[9f^��̢=��)�
K�����`�˖�� ����Ȇ�p	���:����Y��̏z1b��՜���Ũ	��h0�1���a���Ѹk�Ʉ)�µ����k��{�[9fM
���'2��-6� �(ub����Q	��x��99��C��~.7��x�>N�(�`��9��l����Y���WL��ؕ��dQ�~=,N���_(�7��h�$G?5�6�.���eqDm��0���EKf����d��[Ó(u�7�B�f%�$����0ZWw��yP6p�Ó(��6l������̽����'�`��`�\��Q6'���M&_~Ky���9/��22K�����9t�Y&��&�|�uU��7F�E�O���9�\�DeFN����ۛ[)qN. ˟�A(��(e[�Yh��E�&�`����C�u�����"N�@mJ*H�<a�d=����`Vk-�č�s���4��YP�\h���R�d��Ϛ�_�f����C���4!ۺ.��$�y8]��N��W/�d�������麵�n`�y��4�Ŕ:9��h"w������fu�����=���s�3��L�-��sa���hu��C܂��n�+,�/�Jl͒�����mj-����5ۅ����sS�:���Y�M%��N��Yǟj4��uKD��u����08�~SbƆ��I7u`�,�O�7n���~��6�C6�S�+��РY`�l\Nxү�|�"���ށ��\�d�I��8[�i�W��u\�Ky{71��ף,�������3�Tm��\b6�f��i-���}�#�t}ݗ��F�ȩ�����z�g�.<��hX11Uhkq��,��k2��[�b�����?��XF��&�n9-����A�.xQ-�n�g��/�Ka�슗��8Տo41���� ����L�iq�)C�+�L��^��[Ԑ	Oz2nN�ŴQ6`b�>E�D��QSUޞ���8��	�G�tD�&b]��!uCk'�aJ��>����#�]_+lA�s�X��N'D��%�_�0��6���/d`cf&��.b9jJ�21�7�j�3�2S�r��a3-�Ŧʵ����n��I����Vm��/	'7k���m5фR6��m�fy�	H�9b�,ŕ]p܄'9��x�x5f
2͜�b��,K������!&I�(en�L7'������A�<W�Y�f0L���L�΍�{�z���w�5��h�Id#����;d"�ח�����AJN��o~�^��K�L�úlV�ꑑ�&Q�>��B��Y��!]I�,p�j1j*u͠9��I�j�I���h_W4l�\��lb�o�rux�dѣY��3ၔלP���%'<�76n�i���0��iX���As|��d&�����͖��C��;l��9��nK1�}�V-��fA�-p
㫲�l�4b�,�m�օ�#��T��CL�S�	��@	B�'L����q�<M���] �25�i�9��Cf(��f
n��%vÖm��Q�F�9x���R.p���9�T����<��!EM�21�̍0d���݅�M׭��|�j2��p���׹j|�/�g�����[xVq5���i��|^j�w�f��TGF�ʡA�����ݨe� ���_X7�t}u��n�+K�>'�����AY�!L�����c������5z2'~��U]��\Z˓M��C�l���ZV�~ޝjf"}E��>�eb�o�{5���x]�r*:βsf��%Qĺ����i�Ζ-�s�^����{��W�ͅ�.�4N��r�n�k��,=X��Q�w@<8��S���ly���U���妆�1���[ լǊ<�2�@9u�g���IĆLD�s���{�uB�)��V*H�<a�M���kf�6)���tr���y��w�����:ޒu�&<@�t���p���!P�@��V�(3�h��rY�/��Ɂh�.���Lµ(ub6�np���B��E����5�DN��m����[FI$���s����R��+��p6
&����<�"8u�n�,��cfs�4Y'g)�Y>KN7h"������0kc�Mxү�0� ��v�Z뾑�3C&Yw��p�\�NOf7`3I(�Tw�^���+�p?J��'1�;���������F�l6w&ȑ��$�[�՜�����ci�v�,�I���RG�q5hԔ�n��K�I
��K���e�DG�YzKV.j]I~�.�p�˦����i1-�h�$��\�bN��]^ �,��z+�~Y/�e�6j>Gf2n�\�+��I:-�5Zi6�JM�ݿx	�m�Tm�hn�㼽"辭�7W�L����,�5տ�����ٜɗ�X�,�{󫰰.��j�'��X������W�`1p�W�&<u#����3�_��M��t��N
m��J4�cM��G s37q~���h�\�4�&b]��#��p̹��7o�N��c��2#̠�4�S��l��9H�^ղ��¿�AJҷ(u+��q(�~dj�"N�@mJ*H�<a�d��g`�<�!�*g 3jJ�J���!g������u����z��4I���=ݪ݊u<|d��pY�a�,�\Xp�I�۴8��fȄd�u�V�����Z��$ws�9k�
�l}n=�8��o+x���C&�W��ML7f��|�]���B1���ź-�[����Iԝ<k�^�j���,3���Κ-�տ�Ġ!��������p�������X:�z��Z}2r���>n�Xa` 5�ߐ��gu�j*uW�ɾNϬ&�~�:6�x]�,������X��΢VS���R!s���M�S����Bd&b]���3�j-3Ux��ù��se�T���j�.�n����b냡1b�$��/[\nN�˾����25����uz8d6t���Ӥs1���,�P���fe�0�7f>���z.��!��)��v�����&Y@��~��rr<���-�su(�M������E�L�(����,�b:��KX�:�9u�$��jج��^�H��^�fn�uH$��ub�R�.f�q�f��FN��݋��/�e��R���E�7�Ʒ����@sY�pVP����qxlg�#֩9��yc7�~�u�uq��f��Z����*ܻ���Ĕ�Mn��)���{�WຊYw0QGfck�,��"EӾ��FN��g#'Lu�����$]�Tw)Ѭ<��i�v}y.�b.��5e�r�:t��㉲��E:��Q�P�>kv�]e37 ��z�7t����g6���rbҟLfVë��-���qL&L���ت���N��З��Tk���N�L������R�25`εkj���խX�eǩtkn���i�N�s/���Yc1j��[��<�s��	I��&6O{��Gx��y6�_�;��&<u��>P���}�^@W��d������戩u�9�8	�֫s�us!V!�9-�F���&�^���y�IEHj��:��#���{1����V�S�Y�E�H���&D�b����?��s��SI�F�B�&Lu�c�46]4l"�e�O�7\��V�Ȍ�k68H�v�oYf`J��20nƆa7zO2Cԩc#��Kz���N��H����b&�_���f��F31֝�b�9W���58��I��O��Z]5����Hu�8!�(A� ��I�e"���s���f.��Ք�3z#�����3SC�YW�]�qp*y��گ]&�"�j`��K�NHT}\��6���(�D��b���3�n
6��%�����7��{"'i���"f�Z'5hB���"?Tn�y0deQ|S�tw�r�a��;V֘ͺ��Pu˒ͦ��g6'h�Ό����T��_��(~�@���� ���j�։	G]tˢ�-����O/71�^Awo�1l>
à	A�����\����@��mji,"7�*����һiͯ��euԬ�ԉ�u���9T�W5m�2\/2�9��R�f�T٠S��s�9�[���n]W}�������"�g�w1n���
\���x�ͬ��q��8��Խ� g��Jr7Rݸ���eFΦ������䗫�&��{*4���o=���f�X��[Ϋt����l^��9�K�5����~�ڂQS�f`VRͭ���\���L���ٺ��dQ�܀��MC'�ne���b�l�T���u2�ݽN�w��ue֩˶X������&e?͖�݋�Ws����K���7*������.�~xY��0j�N��`�\���
\�x�Œ����r�b6��+�բ�XI!E*;@�,�I������k%�Pĸ��`'�2M�XU0b6u��$]?�׻W��ɂr=�1PM���i*�=�'=#�9�:4G�ɧ��5Ӫ���Y԰�Ufbt�Gn����]GfA?���2�g�{�lj%����u�8!�(A� ��I�oy�����R�q3�/�ͨ)M�p�.�u�Wb-k�]7G�aW��
�n�oXķ"�V���Y�󃍙�2��z�9��,�uDc&<d����q�V�����Nùm�B�	������i�}b*���=Z�WL�}0�	�!�>W��Fp������q�/�C7����ɩ�J֙9��z�+�V�*�Yѱ'aٲ;����s�hB�f�f�6I4E�[�p8N�e���[�쮖11jT� �kٖ�9mo����'���X�Vr��A�.��ƿ�0b*�����fF8�l�n�e]|k��$�,���2�d*������&$e'�\-2su��<�m�r�O�	�l���hY��Ӱ��S3W��h
�NI0'�7I��T�ܜ�E7��ma�u��j�r\�C��J&��d[����ؘ�X���͕_䬽5aJO榞���"��i��u˄�mY4h*ڗ����\rN�$�"��O��Us�J���́�9#6*'�~�6�Ρ����\&w�b����[�uޠ���X��;�.35�p2�EN�sl����`�ȯ�"Pہ�
�/O�d1�>�p��re���۾�吩M�ZN����#��3����+�{�4㮡�k��Ng)����*잪�6C&\un̰9:Ѣ�3u14�����5eK�.��&��N[/��w�u��/@����u�,`��վn��E��k���p�u���;��ru�a�w�LW�:��,�g4��+B����Y�Cfҟ��%�0��Ҿ/f�i��^�/8]��.11u�Z�uX=8j�D��B 3dY&˟LQ#rz7'ӢY�u&sX�:2방��"2�Nγn`�)r!��#�g���^��LUk1��
���ԙ13�]W8b��j܌��L��G��ahToÏ'4g�d��nSw�p��i�_�á6��t�d����p� �R��o�#GN�ң9d/�7/���:;��I����ce���T�ן��$s�S�����L��(u��2�L����`NW�OΙ�LV�(��[�:��æB�*T6���Ġ���B&���
rf�5�1p�joz��p�tҜv�31� 栱Do�4Vt��ag����w@?C͠9��D�S�	��@	B�'L��,o1}�.0�j��Y�Ž�����6�Z�e���X���j�<[�ŃXe��Q/�|�W}��Y���Y�94�����D�.�B�Ĉ	��E{~X�̒��bg��(��	A���<�3�����0��+w����pwY�Cs�L�%dl���ԑ�rY���N&\���.���f���\Mo4���c;��]�h�lZ��)c�P)F�}�J�_l�uڠ����X�5�1r@�y��YBw
���۪�1�z7FML��W��R��b�D�+���z����լ���$_�f�0r�5Ų������K����RX �LC·u�;���K}arc&D�6��Nl�%In�:1��1ܼ�MҺ�N�q'F�ꑩup�i�/`9h�$����MF5l���,^%2`��X4`"��ԛas�W�}rڢS�Z"r�,�0ՑYa+F�cTLA��� sD�̘	AHx�	�vd{��h�,��5j�$ara��տ<l�U6���k�Ţ>� 6I�7��-k5d�6�4�s��8��g�\�+u�*Cɬ�2]�o0'ɯ��4P�FMĺ�~e�k31Ą)�7���։�S};��[h���ke�6�XM�� 7cF�0)�zu��^7׭�J�uDӠ�S�d��po�e�Nk��zǨ�	0p�^Xjr9S�̅b&Ƣ����:��n_d9�~��9����,�\?��11�R����騍ZV��yp7�V��u��̀�BSw�,�<\V��n�R�����	5Wt)�9fRף��nV�����>����YR]�L��1��A51�ZE0��y��uY����"*aJ��i���Ք�!�8����d]0�.��:�97a�[3l��2��n	��Y�W��n*�W��<���˖�
\��Ӝs��m�(�$���
Z6b��Sꖄ��\���8�5p�TF�K���,�]2j������߸Ý��+&����z�6-3�Q���̜X��g�G&�*�8!�(A� ��I�#EL-��:�z�W(��:M�:�VdնGs݀�y��E��Y�k�d�4��2����9=��S��mji=b�!h����27�΍�C�n`m���]�l�s1h�6��f��dh*��,�����&��uO�`g�����͒#'C���șR3f*�o�
�,jb�ot��Y�E��h� �Swb,�ъMX��up�o�^�w�Ó~�&f�u�cj�Ж�����d��a��s�ԺŲ�Ѭ�@'��j�5��T�sM6���!�����fs�~�Y&�{�����As�/��q���_G��ldA�#g���T��G�qx2r��,�S��q9uf��e%���b�Ĕ���ܻFb�Sf��e{.͒��?��r��
C�fW���k3jjݩ�Fd��91��R7`�����i��_h�;��"�Y���4��C���1I,�.k��ٔ����!��cK����ї|��M���,�'i�h�4���C��h�耵���u9=���n�l��0���f�8`Ȩ),fs�����:6pFօhA6�Do�:4�:�9y�$�,�ͅq���4���P3P�&I�)Q�ks���|;k�xE���x�8����LSP�Y�!2W�Ӟ�
��}Y6��MZ�,'1l�(��� ��r�l~��Y&fb�{Z8/w�֑Y���&�,571؉Pw�ɼd�Z�q�=��XW3hj�!��]=�����mA=>.Oĺ�6���7��`�1`��h.4��R��I>��RLI��.ƣ����ʅC���u�PN���>l��Rc�����`�\���c��+Φ��Y�M,L��:8��eBFM!��̚l~%��e����rS鶠���s���wU��:ށj����Y'1j�G�c3���f���0�w�.�q�u�&&}ˮ���V*�ڇ��w)��.���,����Ix����ʣ)�"s���06�B�a��_�+��pաY�K�as���8!�(A� ��I�#NL`��s�>������ X�Xr�ܟ���L	���[���Ɔ�ژ94�5	���Y�l�v1���-H{�-g�����$�+�6^q|J�m�p�4jX^+�`U�G��5<�u���8��A�.���_��6l�)���AJ�իp������Z�Ijݗ㓻9�݈ɖ�eLC���HuC�a���I~�ʹ���1� �H8�J�V��;�d���ēI��Bp޻13�l
���j�+���[l�OTU;n��Rn�8s��ׂM��涒f	�QsD'�֋�dZ6�x0bN��u�!9B��=����$���{p\p�,�s$Y`PL����½�=8j� ��ʬ�EYY35��_�[g��c��_��vԺ��m0g�1`̄)=����t����+��I
��с���>�Kм6Y�.�]2��+q���Km���պ���T蛗�&�l��,�n�%۞�+sh��˺/2���S��`<�`�L4�����Zd�ni,���ⰰWf�Ä�he9��ͯ�i
����$�����9#n&�j��88f����Tw�]8�o�5Q���;��Q���	s 8Lȩ�Z�h.��J�Uj��Sj6^�=�ѬA���ȁs�����~c��c=.���P��P�"���)	IWh�˄���3�|=���Q�$�IrV��Y|m�I�6t���R��(ۜ4�;n���3���]1r���y��|j��\�xm�0�V���`��i��#�j���H20�r+��n"�e�����W����$_?6/<��۪��N�M�)Q�	��@	B�'L�6���0g��c��~��U�M�sʨ1���,k3@���l��7���h{��� a��d!03�Qa?�'�4hN�r��[�d��s��uf�렿���T���G�Y]��	��CM"�
��g��+\�͉~���H~��Y�K�%_����Z7�~����Ħ������.����I��W���]�x��fI�w36-8K��rW�z�6f
�ѰY�+�o&�?4�@�Py�t��
��9h�����x���m*��?2y�@�Dg`��H���C��8��lR�����U5�p͌��e��3F�8�p��c�=Rݦ��9e�@y�P'��zp�Q�x!7��ֹ�L֭��y��\D׭�0m����M���5۽ڧC�nS;UȬ��ƹ5�Ss_����j&��S	���ts����-U7�5�ax��HuQ~����e3��%����ꘑ�&����ج����΂�f�ޓC�.Y5K��OM��6�F�58�V�_�۰��d�$&�����_��ۂ����f	,�n��usc����kݺ-��,�f����9��Y3��Mĺl�*��³L�T�ҟ��L����p9`N^8ǰ��M8�t6f�j�W&��R����g#+�$4�jl�@{�m}z^(HB٢�竹����|s���6���z��,���Z��{!;����%L���bF38�Sa]���$h�uj��/��7ղ�r�6d�roz�p��r:�v���"f�!Y7i��0W�P0O}>��X́Ή���N�uZ�w}œ�Z����u5�a=�V�X�����Ĝ�]�朐s�Xǅ1Nh�r��s2r"�ez�����&<�ɜ��r�hv+�����2����n������#�m���sV�F�»�g��q���fp��f�A���ޝ.����u)�Ni9��[�)��wݡe}�V�ޜ��!s��@�@�Y��b﵎͚��G�&�td�k�n�T���L�<4��d��[��A��~s�Ǟ�"N�@mJ*H�<a��.�0\��9;a���H�6m�	ɨ9�Ŝ���L~�7�f�6�L>4Ps`<Z���J�v2�2�P�;�ϔ�Ŕ��s�-�lnN�k;9j�9�IB��߸�}6cfmn��$��/˗-33n�D�������YnW[N��Wn�d*L��L��â�t؅s��T4E4��ܬ�@3n�Uf�,��s���䯻Ws�=Z8�~���e{���/C�fi.[5ג���]�dn�RS��f��}4wM
��n����a2�hu#p�y�Y�u�YJf]	u+|ů�	K�M��"ԝ-f��¾@�I95u�G����JԺ����Ĥ?D-�S9��:8���e��fb�_T�f�]�p�D�K�.b�,
9jVN8��^���d�-��X��.����\��m'��uQ�7��:��2w(,��VGf�J�b����}XU��Mt���Y�Ѡ1�&snMݘ IY>e��%�֍ײ��̡�\!�&���^�M^74f�$�x�Vg���쟛�΋�TT����@�k7M�R�^������TFf%6�f!T��NE������pb�9Х�"Pہ�
�/O�d1�\���^�������Y0�,�ڴ�󍌚�^����ZV4�$��r�Kr*��������$8�Y�5\0K��)[����-�1Uh�����~�էͫy�J�a&e������Zn�������ȓu�cb�����eŷU_
+���Q�=��uX
nJ9wCL�-n9GϕP�"o�V}��=�+&,�j𖾺g��;�s29�s��9�Є�m3��\&fN�0}T��.f�0<��b<@�9���C�͝��᩻:+�����n�E���ı��R������խ��soz�����-8n�����0é�;�RvJ_�uA#FM295f��j܈)�ùr�%��d���*��vY��.��&ج���%��n^�Drj�d!-���-J�9J�S�Ѕk��l'�W���B:��޵;	ф��Q�Ȍ\C�S&\u�pi�1FνK�y���jvхC�tc�j��]�C�rY�/���@F͡���d�3�ͅyƘ	�����S_�0qh�_��Z��Z�ӟ׷N�BJ�Ry=���>�T��ȬĪ�s��$9�.�^�C�4�\���u�8!�(A� ��I�ï�>�pYk�ƍ����s��!S�6u��Q�rۯp2f�����,1j&������2�f�s]��^��;�.��&Lu�z�S�)�Zd�� C&Q��5�$6〜�G�f=�>1)$E�[P�f̜5b�T4�9��|��Q�~A9�V����owY�'��L�`8������9�.�d�}X׳��
�j��ݐY���o90�ʮ4��D-1!H����Y'9gs۽��s#�a&�Z��趓Yg�C�4a��(uK���_�"����ۤ�̩�fs]wNn���N�͜��tZ�J��沨�sȎ�;���<IM�s�V6�̒�E�;I�I4�u3I\/�3� ,��:T�>��uY-�8�߂����9�Ѭ^�?�W�Q�fa\|ɺ�,�k�f�6:�����#3��y��0<J]t���:�Y�K&LȊR��b6vkG������MT�(����0|i�}n�aI���"3�
_�$̈́���-g�Kn���u�f]Ͻ�x	F/�n.85R���|6��fo\6��#�����P��^ͦհ9�N�0�mf��8/��c1�[
&C���9��&��h��_19ǫ��G��vn�h�7�i͠3:��ek��͑�Vv�3�p��ȉ��B:��rX��21��bNN1I¬�������M�#�Ea�0!�X7\�\L9ko��d	�[�26�s&Ą ���Y�A1j.ySik4+��۬����Y��l\P�����[����SrS�f�j�y��Y��tʒ[��Ѭ�]��*�>@�YtY2��C{5+��k�������"Lu���١�B��/J��ZW5'����~�_nd6�L�h�d$�"���9���\�X���dOש�9�g9WX�1�����h6���[ML���s�@��{�9�z61�^�U�f4��;H?>�c&�^ ��������W�I�_΁��X���;�М^`�n�ĸR<�jm��5 {��lr��ɿ���m(r]ʹ��E�M�0�_
�8�'cq3�cA��q��?�9j�ci�m�f��SFF�8�ݽ#�t;B�]s���*=��,��+�M�[6�qP�sTĔ�Y��(�)�{a_ �81�l�Af`������df���� }Y�9��4}�Kh%w͘Iʺ��uyP8��\|����&�72�y��a�N'D��%�_�0��d�W`��s�L^1Yrcpm��j.x��[`̬e��:/LC��ee�2��D�9x���b؄����(�$�����in�U��E~ލ��;��fw�&}sӸ\�U�6h\�p��ed��>d��1����)�y��#�d��-f�����8b]�����̍���G��3��M5^΂�f�<[�����VN�!u��B�R�FL�H̐ ���,�	��.�]w�_��B#'	O���p�]4���!j��\�5Nbh}�<ƹtnE�K9�|刹�YaaJ�fIɹP�"j���c!��&Y'�9p+�<^��^�Ŵ�r��B%���
�+�٬��A|L�5ژ����ud��8B?��_��M�W.��1�Z�erzm	�&��Z���=iղ]�G��4��~��)51�<o��SILĺ�8��um�	Sz1j��xG*�V�z�S4c^����l2��������M�c�	���"��)����Z&n^h&�ЛY��+��b�D�KiY��Z�s+<������[��
��r�7�1д�w��aC�����@65IR-2�BFLe�}X_34��D�U\>r�l�����y¯�v�7E���� T�~y�$�AYL`���s��`��|��Ԧ���f�o����]�\�bX.`6�Z�����ͯ��5	�jF��{"e��Zr��Su���1M-�����v�`&I4kxܬ�SUy��
]�ksC�$�z<��Ӵ��D�+��"��&�,Z3b~�ܐY�˂Lu{K9'�F�İ`]�f���j�������r���DS�6�3����L��f���&W/�޲[�׆��0�3�
Mx��a�`�YG7���&n�`��IQ���qh��(HQ�����l7KR�5X~j��bܘ	�:2��!���-Bݑ�D6��/�bb8����`��Tj.�â9�v~$�o��f�V�ME#�U]�7����[`�i�X��mQt+/'L�Ѽ�õ2Yx���m�uI�G�{J5b�ʥ����� ��f�_�}4!RGf�J�b�[��3`�A�&���.簲�հ1�9w6m�P�r8�Z�zatS�~�Yhݬ)5�����Y*K~�ԄGh�xV� '<�Zו_���f�����a��Ʀ� �9��<L��Ȭ��fѫIr(J]t>_��ku̘Y?7a��"N�@mJ*H�<a�d�����戾���5�IΦ7�f��,����l��b�����o��p��c�����e��}6k�F����ܜN+��ƬQ�n�nH��8�n����q�+�ԭ̓/_7�[v�
_!k���L����<eN�ը�/�Ux��/f8�:5f�uS�7��nV~��uԺ�ލ���V6��T���eݔ�d�;+�d� :�fW\��/����ʶ�B�G5L�m�U�43�L�j��{ɁiYW�%�L��Qe��uKu��P�9"�T;��Axҫy۲��氥��_�{�f�4�䈚5Yv���^�-����:��_.1��m~bm�Lש9�?�S ��ɷ�Kjy���=1�u^h䐉1~9��4��	��ۑ�4�11��Yӫt/f�{���'�qC�P�p�l}�x�lt}b�h�fYl��Mĺ��"`shY��&<��fV�͒�#��-�Su�A�L�ɋ��p���ʀD�������4t/T`�,2�I���g��L�ld�͸�S��pD怼&1~��=;76m���uY�M,���F�,�]�$ҳ�M������碬u�8!�(A� ��I�5�h`�\�C���j�u�6��4=�wꠑ3T0S��Y��Y��~r:��.'8�.k4rvG�[1j��[5I�^�hojЌ�n����m�}���	h�Y�[r�/�Q�J����2h3�
ŧ�Vr��*<u+��X0?�$����e:T_3r��լ�4h��o�J5�4J�I>-'�YG��-�5Zv��5�$̺-�	f�pȨ�XW�_��{�hج4aJ���Q�R3f5��Y�5��92r�$����t��s&����y��*5p
���_��W�t?J]�rn[��g��a3�5�&<pu��YP�L�aH��{���RS�=�1�F�vp�l_Y��l#�5���S�z�9�����A¿uۮ�f�y���!� d]�F�C����g�Տ�߂,�͉�:�n&b]����C���%}���X�h�S�qBj;P�PA��	�, +|�0�f).��^w0C�nZ�+yXY�h6p00S��Y�6�ny�) gy����FN�]�Ճ�J�㸯�^g��_%9QӋ)u�a�8j]���Cܚ./5)��u��"4j�!1U�u8΢��#&Y���u3�]�nȜ���`���{i�Acf@���e���_4+q�>�%ݗs�ŘY��6��Ѷ
d�WM��K��&��m�T����̡ N2��l�E�z�����2rԜ�6)�_g�~�X��f�`Fu6f�p,B��t������9:������9dn*�huf���Ŷ�Eb�A*�ik��#��0ՁYO7��)�&b]���ld��q�º�n��Ymf��I�������F�4�7��:<�H&\u+��#�T���u#5��� ���䂽|����(朙�S#���)��v�����&Y@М{sT���}XZ��VS���
q���¿��w����l.�g	�	�.�e�P���R�8�����[��(Ƙ	E���.���Yg5H�l
��l0dnE�[+h�Y�%�&i��"���9.ȄH����z�19h�H9���s{V�Թ�ܬ��I"e��a�f��x����W3+)�L��74k����g��;��;<��ʁi���t�<�o�b!��ۘ���j�9�wz2�WsC�J'�4R�����g;1IrG�[��v=6A�O��|ր��9a+��l�0��� ƺ��͏٪�М�bN���ock�f%�"��y@rsR%�G�\�u6�.��������&<�7rJ�3�T9��������I֝w@�FN����7��f��d2�ʱacf���v�ߋ��|�5H�o٫98��5_�+������X��٬�꘩#�f�oӧo���uY�l�T��`�e/g��&F��qެ�:��X����f�]�x/O��f �̸Q��Y�,��.,ug��U3�6	�����2=b�v�Z��4�Eù��<��_�$��E򲭖�8��4�w�Z)1aJ��o���9���&ܰY�`V��j�Y7�v�W�lP�&�j��$��n]�<����!S�qBj;P�PA��	�, �<� ������ �5�IΦG�S{G���c4Y*k���w����rD��:J���W��o^���a`Ԑ1sլ2a�$4\�l�r[(|5l�B�g�]v+��'nx�?8����q����^ja�&�q��C�f6�2	�"չ�L�vf�����fԮpdfVf	�QsA�I~c�,����%�l{�����Wu�x���u���$�iS�LXҿn���t\dj��_�q�fq�I�s$��Y!b�4�3�͐��?����b������[-0j��G�c3jlry-�$����t�{ˡ���l��[���:���WÆ��u�sr6����/r��Q6��$���917O�M���KΡl��7$��� r`\�Ei&����1s~�i�ŀ�Y백�C��6�y���uYx뷬�mc�&��_��_O3h�S�qBj;P�PA��	�, p�q?�<���B͜['�٨�4����n푁���h����s��d��>���E���ć�f��!R���A��^ �!%T4�b�Ą�n��1罜0��:3��!m��&I�(�E���/3bB�od�"��bY�d��c;�u]6j�l�Lj���2+���Jl*�.~2+�P�9�c���>�1|N�E��
J 羑Y�d�L���a�V�b�M�IV�ˢ[<�l|�j�����b̤�\w6��-O9d"���so�f�OY1�I/͌V�W���xF4	�_78`Vq}؈QS�Y>b�|y��0ՁY\�w��F��^��3l%���%鶘���SfL��^Q41*�9k6��0Q�o�MF�7g!4l؄'�0�
g���7rj��_�k9V�Ir�S�꺁S]_��5[Ǎ�#�74b�u¿���}��'��Z���Y�ŵ���+���6yX�q}�����D8ſ#�x*&��5;���9��4�尼��џ���^%4�5m�[�}Y�e����-�s�@	g�D�˄]H��F��*{ҿlLv3�T�{j^3h��L1��$�i����]�f�$SG�#sΫ�9`����_�x�_&�h��]&����tK2�BM�o�^~bĬ,�C��uY%0�S�i4p��0�?�6�\70b*����υ�`FM�S�	��@	B�'L��,�����|VcI-b�é��4�ٴ��K�xj�)hAcf��9���f:��)�.k4r�G�3��?s�prL�YJrP�2ၔ�Уa3��݄D�,��e�es�
O�������B���hA�3t
Oݡ͋����V�:7��s)��I�?�ȨA#碪Y.�25�c�x��I�zg��t�Uq�l���.^3I�n�J�YU6r"���0�.2ſ���vY��\�߹#}!<!�$�"��M�'���͐����uXX���"ShNj1�P�t?J�Q�R��8��;X�9�,�Uu#'<pFf@� ��b�i��|XXN�"����3ae�u�T�7�i8���S�z�9ԭܽ3��^�:1j�m�Y�fb�����������7r�c��E[�C���uYh`���,Z1�I��Kp�Yύ�!��)��v�����&Y@�~�0�y�����P���#�p��8��)0��6���+�Mj8��uP�FN�]8O�(ǵ���0�md=�$�15��Z��l��R�u������"e��.x0���)�*��l�,Z[9b�u˖��ޗ�!ki�mb�Kឆ�n3�|4K�x�#&a]����>�АI�W3��}21]Gۖ��ʢI����K���l�Y3�ƒɷ^Nֲ\F�n�娹":6)�_w�^H��|Ӯ��9dFm6f��#p,B��t����[4���l����Z4��%'&�hu[D�Y�p�4�:1�B�F�U��&<u�"g��;���X��_���l�\�Yw̺�Y�Ѩq�޺�y�����������9Wα�ɉ��:1j���� ��X'��j��̠�Q�Rw`y��g)��.<E���� T�~y�$�so�
��a�]�O�%Q��lz#n�,�e��ko��fs�Z��r�V ����.Y1�!P�P���V�(3�h�e���_r*ЀYh�E2kL&�Z��%���,��[�j���q��7�fyW���%pH\�;&MI���;��w�s3��Y2}Id�j>O�*���Z��IyuШY��f�7D&b]6^�0k�6��%�{�͊�y��r��\,du����ʺYw6h��بin,E3I(�T��uD��NL���Ĩ�z���s���������s�rr1pb��Gs�����b.�S{��$�2s��t��|��������I��Vb#�~�n"�e�m���Y���%���5�S3h��n�7f�@#'Q��/6� g��S��,2j���I&_����݋�FN��"3��19I���Mq�[]wߖ�;܈��
�Ѻ|������,��/��G�x]��nAd���<��#�6���r��X��|2�qs�Ws�Ó~)�Y�eq��T��}+x�>Մ�n�!s��&A4Rݶ�8˔��NZ���,��P��Q3��_�$�V��;��`���e��\hl��@Mxҟ�l�l�*��e`�@s���1U�&�f��r�*9����s�du���g��ݦ7I��)��v�����&Y@�{y���0�=M�4`oFMi���z���d3�d�n�����.�Y&p�=��G��-��[5f��΁y3�p@ʒ�s�<���sW�"�~���WRL���Sp�u���8^�7���"�q��#͋��C&�_�:7��$�	�}1h�lέޢ�y���K���:8�k��n�t�5q����� =�Qo�,�E�9�
�!����e����j�k3��MM���%��-'	Α�4��!e�W�͐��?k�L�B�&S!GsR�5I��Ա5��9�%i����/�u��/­���ۘ�ܩO�pg�܈�XW87|��/r��Z��ܕ�8�}6�5������P��#�L{�2�nY_=31�_�lȘYrl�Ԣ�a�u;۞3��uus��>4n"�e���tI؈	G�h|^j��~��u�8!�(A� ��I8à��"�3�f���RS���qHC����]2l���,�f���Yއޓ�C�ٜ!g��-�l��H݂#�f.6�uH	Ϳ�:1a�[��\�Y�o��[���lZ�;��~��(�2#&���B������,�
��Y׍�Q�p��v��4z�B�Fκ�� ����6h�,�̯���l�sL��s�n�N����,8���
�+~���v�d&Q�f�K{��Z�/�1�W�1�1:eq35�B3�����\`Ȅ'��-�a��9�Ժǽ�nФ00U�{7ѹ��l�J���]�-s8��:���`��-�3n%���'��7�u]�Рi����ʋÍ��2��a���&b]�Oͦ�L�A�7�I�f��%�85��/�{}K�$9�f�_��T��-�=O��>71����nV�(o�����88�I������A��+ݬ��d�Y��kc�� s�YK���l~YmTL����S e]�nVd�o���B��j�ǑfIv�cn^ΑD�ML�Ý7`ࠁ#�LĺL���8��*��G���8}W����g��hbR���,�u:纊���Pw#1�#�=֦�l~����I��W�r�L��M�~A_�
�c2��Fjb|[pWi�7r<�1�.�ys7n;8�L�ғ���Q���]"r�Lm�S�	��@	B�'L����F� ���.1`�1���fԔ&9�>�OE4r�Zfj��
�,0@\LS�e�FN��(u�/F���U�����:��J�9G��A��Nx@�i��c�W��[o���o+Z�{ެ����,O��^��?�$�����:�\
3r�����9��ek���z�kN&Q'��������6��X6�n�3$�[7r�\�E�&bYq�TZ<wE9ŷ����b��(S]_4G�
8�$��m۵��1�Ĥ�_k4�q"'S4'�R�&�~�:6��E��8c�vϖ��\nĄ�N���p~d�.��U^�b��"��6��Ȍ��}6l.8��#0Lu�%g����0��/B�2\�Ew3�-��'��:r�^/̒D�p�\����>�����.o�r1��9d>����XO3h�S�qBj;P�PA��	�, �p�0D1G�1�^w0C�nZq39ܬ��f&�.��f0ˇ���p��boؕ�m_w8�`�0����	O��b��Ep�DM/��-��BA���q0���� ^0)���Les7�M�T�.�
�J7 Y��.���MCڦ��癚0խ�@�:��IX�n�Ű9D�ѐIZwv���u\^`*�N�͑�_Y41ƿ}��J4l�Ƣ�2�m &�a�!i!h?��5:��S2��g�qͥ�)�CfTfc&�:
�"ԁ�N��:1��R_i0+I� y��<�!Q����խ 9�C0� ���,��9]W5�T�.���b�D���/;5� �Y�t��s�_�Ѩq�To͟n�6����ujԬ庣YJK.\u[���mvCr���R'f2���n5)�u�uD����({.c3e���A&BS�	�� T�~y�$�J���s��ۮ��S�4�YY!/��3����4.Rx�tS+r����	�����_��(F�	E��,��|������^2�y`�$܊P��q{�٘���+`MVc)�Y�
p!P����f��4Id���E9�DM�s3�Y�� �D3G/4븨��t�8��0�$�y��oxu՘�XW�[�\�#z�Ԅ'��G,���;����f�$���q7��EM�_�بiޫY�$TF�s�'s��<H��(uw���XZ'J���D�U�4�l��9,fng���^$��r��]�f��l���O�w?��a�2�[��%��N���6��.�����X�Iv<��s��9�~�t;��!����f��,09ɺ�o=�ć���)�`���a��T��r����y��l�~�z����l�/�e���Í��V���}e�,��̀��g'C�%�f�"�c�&���oc�A�ȾLn�H!GNĺ��ͬ����Ԁ��fV���)� �M��no�S<e����l��(el��6q��I
�UsZW6��fZ��D�vI���s�C�9�#�eᬯ���8�0�_�W��BnM��L�|`\��21`М�+vz�Er֛�f/���I��l����C��)��v�����&Y@�{y��0C70���ͨ)Mr6��C��@���`^�����Mp3�
ζ�MR�(u�/f��k��L6��͂Q�f�\k6f���� Kn]��a�FNX@�u� 1+rk�EN������T̋�/�p���w���^�2	�"չ�\�vf��}�0��=�4��Qs�.��_�d���ӓ͆��N�Mݺ#7�Q��-�l�<]Ĳ�5��2���[����Rx���n6��_��l���I�_$���j���Lr3$-�pWo���jd�Á��$��j��G�c3*�a�F�ƒ�c�� WÌ�
�2ww)�Ir��6�p+} %�.S��C�D��MV��d��3�04��q9��#.Lu�5\X95+�_���z������!��= �fH�|_�N�uX��G/9d̠�� eNĺ,43��L�z��Q����w���CL�S�	��@	B�'L����� ��mAc�T3p6��3�����p�L���
?�9�V����\�C�\l>/��VU���#si��_��$	���21�([8��.��,'L~���8��)5�$I��E+��3bB�/h�Ա�f}N�e��F���f�����u=�����U ;AV����&���ܬ����*ԝXk����obܰY�xw�T���M�k6�d&Ywp_1l�ƍ����a�\��s�f��:�T؏PWܿ�b.�����H���9�������	g��(݈AS�a�Vr�����b9��K5L��%r���qz�$��6�f)��m0��*�v��Iu�l�t1�4�j�͛�r��I���Q�������s���f��Y��hSj���[.|Ko��/�����,��6!W���u8����e�i�lzȜf�71T=q����Se73x[VhȈ�3|��1sxZ�3��|a[�e~2%e?)��#l�L�m��)��DcSw�>9�2b"�e��9��AG�0�ws(:?��_�;T,Hψ&&���5x~1M���f���bRG�[��,�����
O�-W�r�L�mvu��RsI*�nO�e�&η�]8۬��/&b]泜tpV�1aJ�,��͹��2���9��QS�qBj;P�PA��	�, ��.WS�1g�B�ʫ�5�i�8aO��}�c�����x8`sK:��.����9	��ԭ��|��a3	f�#ǐ�S���@��đw>�2<  �͹�(2g_x��/�5pnDE�i���
g��:2�͋6�'&I�Hun.�!�9��k�f��V��Z5�6����r�$��ȑs���n	.��3s�1�$��LF6�7T�XW�?��l���)�EN��rD���Lȩ�o�H^�'��D]$��A�����Yn��%��-�58�7���VhN�3NM��(ul��#x�bb�wn�ۙ��FNx����U�g&�!s���Y�E��-r���z��|e��n�D��#0Lu�%�+�F�3I�E��f������!�&_4O`�fM�l�i�&�n����{a�Mĺl��M�A���ʐ	O�(|>
��
B3��Z��"Pہ�
�/O�dY�a�0\��"3��|�s��)M�2;d-�h6p�6S`v9��g�IQ�v�[��pԸ��m��_��\*K�26uf����Q�NL�[jh�.�͠�sk��S���u�8d��Ù�*�ʬ�Y��r�$����'wC�M����S�9�P.f1G61	�"խ�6��e��L2=�f��C�����k 8+�&��嵻��s�0;��._8�� 5r،��l��6%�v(9�'��f��Mc��73g/�n2}�E��~�ub��b�'GΉ¦ y���w�Ť@�na�i�s���\�xVs�_�e���|���CFLĺl���f N����{V��71�$\��^Y���k�����&V�ͩ,'���eKό5��� ��X��p���2��'֙9H�	��qB� ���* \l[8�,���&4���u��d����)Z] �!PG���T�3��5�Ԁ�?O��dN�C���5&�p!J�v+ΦWnI�Ij��+���6s `"u[�?���ņ&�h2����[^�܌eKkS}��}oˉ�� ך#�]s3I<>�Ő���,1��+x�-�mW����?Ժ��eX�K���z��b!���s�����N�[57���$�E�s0�7l�l'&�~����+������o)��C3�`C榮�ꈁc�i�f�:�Z��\Ŝ�+&��B�lРY;3�Uc���ݸ�N�v��	n��ՌX�Y~��V�6�%��hC�rjԘ1S�^�&f�/�h�$��X�C5z�]l��9���,˛	�p��57���Ts���^�se���T^6+h���n��YtC��Ae�jjr4NK�tL
��
G���ǲcׁy�e/g����z�Yot�.��N���aJ/G�v�s5p�+Ȫ��హpԨ	O�v�Dl��Hu۞�pΝ��Lj��es��t��fx��c�������O&b]���1W������u=��6hN�g�)[���px����`繛$ˣԭ�f������Z��"Pہ�
�/O�d9�������8p#�3jJ��Mo��{�C43�[/.1�����?��uw�&�u���?��ߨ3	��By�.6��p@.���^e5�B�"�纺�s���ӻ9��a��eঢk���C��Ԥ��VGf�@��7H�����Z��3�d�ݿXb�,��-��cUͦ�,��L��@^{�u�\603�OAjԻ���@mW�_Wܿ0�D�9ſ����Y���ubSq�f�|T9lԐ���H�s���]���Yn��%�掹���2������&A�HulF�E�ѥC��p�>�6f
H-�f��e7k��܋�lL���&bYV��_�Ewc��p�,3'ϵRSY��{	�q@�M����HX�j��3I�E�;���W�L�7�º.�A�}F�p�\�8�mJ4�c�Ѱ�X��_���u�,�Z�z��bj�"N�@mJ*H�<a��0��g_��¹��u3�}#�2K�p�L��u���i�i�^2���8):t������A��q"u�d��Y��0��������9D,�LN����n I̙�&I�(�E���/3nB�o+�$��7m���4q�u��I6pАɢG�Ss�=@-��u��C�r���V7a�[�ŵ6��Cp�:1�nY�Y����*缞�C��V��MH֙9�-���"i�ۦЌ�c#'LuM���uJ���*, �97)�N�;l���s ͔��ɿgu�dY�w�_�fэ�ĭ[�̀����S���n���䫾�|�9��k�f���uK�<^����l�����:7���%L�Zpn�z-0�`�����&RH�mؐ��`԰1S�6u���c�J���97��]���b��fb�z�}��T�V�Z���9듾��8���x�Â���&4�}ت�<|m�Z�������d�M[K�̍�nߔ���|]0r���y�Ԭ�?�~_�mWr#�[n�O�Y��U<[�0�r�U]��>2QS��,V1�{���c]���Qg�]2`܄�N��3��=�#�ey����犩aSӻy�u>a��dz5bΑۼHД��eKK�1��f�2/�C5٬�5Z�5x���"�݇M��z3I���m�N+�	6rؘI�Ws�_���L%��A�Q���b܇sO��u�X�G�S�	��@	B�'L�����>�pY��V�Z��DbƗ����~#x}��L���q�ܨ�F%󂵮l�ǵK�y��r� ���	�28[�9������(~E��d���3H�)XW4[M�*��.�ِ͐���뾴ĨY�7t�`Sٺ��?p���:hb�Ԝ;�x\��\a�L7�HlR���A�<Ĭ��2uj.�C�p�'Y��r�|��7��uٿE��������	S�7-`�Lqq��ߓ���c��N8l�v騩Ư��s�����w�F�Y�Wx�'����Ac&��@�`k�����l`�4o�1���r'*����w)�I��o����Z��uſ���]�TLx�/�d6F̲�}d*��؈�Nk�&LuO����hR�G�[56l�+�@�I�7s�-�z1���fY�?3r��[�p��j�օ?ur�lf�y�;���x37v���e�{�p�q�'<��� mb��׮/<j�r�M�cr��!�3U��0�B\�j�Tw@U�:�97�G�[_2��ԅ3HI�_қ��WM���7q�����q�v s�]rd"�e����͒_`��	O���j�q3h��ώQ�0�j1V�u�|_P�,���EQ���$������]1�T��ê1M��b�6���\��;X&�md�}A]�J�'�X��AN�pVa��ַUE�˾��t�.o4aJ�^`�౱(���b���ݦ�$��� ��,�u;���;B����y�!U��b�\��f��հ)�:T-^9����fax0Q��;����؊�>
�V��������N'D��%�_�0�b�m}��r.,'�1ۮ�	��4�5qsy��hֲ7#�[o5`n<�
B`�ͺ�9��$lg����l�	S��W~E�,�*�y�/�w���0j}���]�;P�v�f���T�l������SeZ����\�$�6��oGe����Q7r��2�$3���.�ӌ��[\W|�W�L����,m4�+PNH#�m�D�lnQ/�$���F�ٷ�Mׁ9�����&��u;ǎ���8�P��r.��wASz6��=7�C���F�^׳[M�n�y��ru_�Ѿ��͡!��j�\�f��ygU�ͺ�y�5�A����,�s���~5�G2����އ̱o��Kg	����<�}8c���W#���J�����|� ��彔�����X�rl	� S	=��Z�������ZEgH����~��#La�i� ����lxxP>��A�p=R������t�&麙����i�݌�bVnh�un��y�����e�O��=L�I�h9�.�"A�Tv�½,�ŀe�V��]�bB8k�	9g��a&�C�p�9�/5p�ʧ�Q��ص�3����:��u�8!�(A� ��I���`����\�QΚ�bi��鍸�Qh6�x����oģ�9���JQ�V�%:ޖ1�:2f�1����+궻x�"��񝬻tg�-=�+���1�z\G91s��D3�o���|�*�73f���:8�~!o�71�R��p|�ȁ3�O��z�y��
�ax1/Z4k�6Ij��Ѳ�rpZh�7��'�Mr�m|\0�TFG�{F_�Pc4�;|hZ(���nXX��|&s؀#�nuh�kc6���Sw$�O��V�#ԉ)uh���e�o��N��8���	ɺ*����n~�ߚ�9uאMJ��u5�u��S��Q�����3�d�%t�/��]-8���������e��A���!]��ݭ[�6�׺��6[��&_���ͺ�rb��YVp��yT�r���k�����t�^lj��[C1'01j��뫶p6��ŗ��%�t�pg!8�)�/�r�|�S�Z��׍����άU&���m@�=s�o�������M�w����lpԄK�ހ/��0��RX��w]�l�n-�sr/:6�:6�S3fo��y�p���k�B�uG���n�)B���l��Y�8>���F��ڣ)B���cd?a��i9h�D++��`$�C�Q���pԽ�1?�U��؜�rܜCjĄ�nz�Sy��A�.�lfT���tM�f}ɜ�{b�I�_��<�YI9��{��$Ǎ�dz1C�uZݮ[*b���M
+R�}8��0��/J�=t3&��fb�ۼ��?����Yv��p��e#s0Y3p�D��#�)��v�����&Y@� �.`.X1Or���F�n��h����t�w����'��moԺ��d^�֕�!l�R2��"�P�Y�Űqep�N�q��%	Q��V�1!g���c��0æ������5t�u��h���9�l�
t�V��jF��J֭����^�2��2]��MJ�u_�`�P������3��FL5�'Y���ܷuX�XW�[�+pY�9,M��?,񃣛�Z�?���lvy$��&C��^�ڿy�,�d�\�d�a� j��T���!vu�Ձ+�~�޺�m�SA�hsn�S ���5<�p4����$����I2oZw9p"�e���R��2j~sKpW��NA׳-��G��0�=�
�?��$��n�N��u��Ťu�9g���Ӳ�f�$�wl���>W��[oj��Ȑ��[�庝��
FMĺ���ey����	O��ri�llԨ�����V� r���F�C��e�(ĸ�Sջ�fN�M�Q�:27	�u��I�R��dϩgz��&͘�m��w�s�>݆$�m���~�6�R���k)�A�Lxү+���9�-]w�_`6�&�r6���\&�E��̓���>L�Ys1������T��do@#̓���Xl]���|�i��M���%�\Ű�uK��w1lLN�pV��[	7��*�$g�rN����'����Ɩ�BptTݻC�7k��r���;h��!,�_�:5��u��Y���Zn6�x��9M�`-b���`ؠQ3�T�.k�fجܺo����Q8��j���s��:E���� T�~y�$�����ˡP��af�n{�K�Y�7Þ�������u]�K ��
2ۯﺳ9��$l?/ɐy��CS�����#����=�����$IvS�l~��f��n�P]�Co�l�����*צ�Y��t�UY��%����|�Ё5I�%�(���Uשas�Q�kҿHuh:4�f6��HuD5G�"�t�U������ᰩ��6cf�o��8��� �c&bY�m���nn.��u9�����)���/[^'u�N�fWa�WLNq}:��;h1�^(o�0�LQ�̃s͠�A���a7�p����9�<���o�&O�Å�N����]?��&�~۲Bs�y��[�-��ƶa�5G6��ҍQ�.�Ԣs�nh���ӣ�����������=9��UQ�.k,��¨���+P�1G&)�He��nþ4	�#չ9�_44I��H��:���܌�ktX�]�25pn.��PZn7�pS@1d̨I��̫�J9N8k�fY.��a���9)�4����.�fb8$�@rD�����f�����M������M�:E���� T�~y�$k�/0� ��X+�
��'�Y��lz#�����h��,8�M�s'<ԉR��KpU�G��D�.6k� $ĄF�u����#�2G����!���edfc벎r����kx��nX�8��!,I1hμ���Rg.�����06J�b?�7����/��p�a�\��ڑi��M�	��V&]��շ���~��}2n�$!�$=�����Mt>Ga�A$�+νZjР9�P.G�Ss,m�9�u��3#�,[�d��S�*��݅�N�:1��p���5ۿ씽	ɺ�t 9 /�*:��{�S���ԊZw
,�x@�t?R�U8?���K&�p��{FN%�q�g��,���o����lA_��n�zkR-2���6s:ɩ��v��Y��BNL���%������f���_�Wg�v��ԉ� V��͊9��I���j��:�aS	s�^*��;�L���da;�����������ḹ��-�s���fb�����o���ݸل�3!�_3K�~��w <�Yו�����9�S���x�A˫Z���sp�� �:1C�M�YɊ�-����
�'a��r���c�\��V}�5�ؚ�I�z�]�oC�M��<�����¹����#D�ʉ���TU�j�	C�����'F���̰�xS��G̭9���τ�#�M#�.�.L8d6��&���P̘�pJ�	�5_1��l����\�mn��s�8�Twu��f��E�[�g�B ��Bl&ƺ廄6�zj*	�eg��9�%�G�����4����He�8!�(A� ��I���.`��y�.���F�nZ��kF��x}��L�T�,�czYmMN2yf�����Ჹ���� � "epV�_�e~_��ůhu��r-I6�Yl��9Ⱥ����,[2k�&%��1�͡kɟ������.3r6�&Yw;o�uVC�pc����qؤD|������mL�vr�Kz��Rɺ��.�)d"�e�nǲZp^�N���։�J,z0�G1��.1b�F_0C�M/����۲�`�f"�At��\8����!n�����W�r��yx8n�Z 7u^q)@�Jr�J��*����Y4I��<���Yw9ˊ_��ff�o|?<�/��(�X�n�T4,�-՜���0�=�¹"�I"3Jݪ-̃��_ �$�ߵQN��b8�#�$�p���,�c��cr�\�es��!W�}'�"��&b]���r��\�E��+w�y����i����3��&ɱ�\�9����S�[�kg�Q���ik4�@�IBK���%�xNݥ*�L�p��88�i��\3w����Y�單?7�R@!�TѬ���u�&<��B���9y+�㺯�0��̡ͺ�� {6m�͑��-m1�e+HͦmkQ9v��Y�3{��	���m�4Z�h���0i8��e�Ƴy}�mM���E�=9I�ߪ�+RI�.���C�G8`�)�8�L̦��Ks���n)� R|�9{��!�.���_�Ԭ�����fi�A���i���[�8����kc�&j]���ϕm�q�N���8�F�9��5S���"Pہ�
�/O�d1�>�pf�B0�!��P�J�Y�Xw��{82S��"�us'#N�ͭﺳ9��$lgs.�R`��a�[�lVQ�S�@�\Vs\/��f�$�������t��0@Df�([��Y��lаAS�Z58l�qEŨI��5_�Z�����L�廄���$Y�b.�E�j�_��͕?�Tb��R�|VȠ��J%�2R�B0�3� �dո�F� �1M�e�~7q�-����	r�E���-9f�j55aJ/�8CsnD��>7r^vPP��;����^�lֱ�w��9l��:ư��9�L�W2E�뼹cM���3c�
L����4�j9f����{n�����X�n��K[LR�%���{���j�\ϑ�`��u��f � �Mĺ�s⹱~�RNx�/�MݢW.�d����a��9ɺc�#��q��뻩���I�E*;�����h�G�ss�Xjh�P%ӳ9����'�Bs3�7����g�.<��V��#q�_3j��=�x Y&n*X-�Whu����<x�e-��}�N$9C�ՌAؓ-A2d��M-[��8[�8�W�y��#f�:E���� T�~y�$����0c�j\ڛr�Z��$g�qs��\׵7S����A�q�F�6�y��l���s�/���p$�P}��ō��Qd�l���M�e����e���,�p��VRL���κ'�>J���@�|�uxү��8�_`IH"s����P�Dj4��ŷ�����͒9$�糘���Q�L�3��4ၤͭ�";z����\�/�sb%=��[!i+7}�9��Sw����A��N��n����z�5�s�w�%5h�T���Bz�p�����	&�m��Kd������9/V�Hus�ؿjqv�z-C20|s��sb#K�}s3�6��!#w���%����0I�(u�i7�&3h�қy�K��tn��9G��P�$�B6��sm���z�9#6�B��#�H�pn��6~�� �Y|������EG���>D�+։Y���9c�T�GO�~hV�E㦀��Kh�jqɺ��[�#L�#s�d��Ynh�S��7h^|o�$Y��3�Ut��~@u����ߡh�_�{b�%UmTRCF��,P�Ы��2+a&	�6���E�C�I
��C/$l�_8j*b��b�n{��ta�m+��Mĺ���Q��fܜ�r��]�p�����&��J��ԙQ��g��)l"�mO�*ZF�D�M��5�E1]�P^F9�dЬc��ZΓ�Dp�D�����_��>
��,�[��W�L��r��k_�%��'���Ί�'䒁�&��k��nh̐�SiO��uC�+��M��Md�D�K���`�ľ��u)��a!�ݰ)��6C2q��-ss�ZE9g�%�%J��Wc�IL����Υ��ItW��t�c�*�sJ\��u	ֲ�-��q��Q8s���"�E��R��"Pہ�
�/O�d1�H��rO�<���&��jJӊ/w7�bq��*h�r����7�.�P�Ysjl~�7��[_l�Vw�\��nuh�u���$O����f�6�Ĕ�u=8���h�T�T��/s�.�d�M��c�����A��q�ؤd�X���?���Y����]�22nԤ���E�Nh�ΒSY��d���i�,;C���v:5���C�½z���_�s�L��s��0��d�C��{/Gͷ�����⤐𺛽���U�unց�b=��0�-+3r��!Vם��esw*��z��5ڐ���2Z�ai~�S�_�u�W��+/f�`&�72h���%�����*-}7n�� ��o��y/��%4���
?A	p��A&�^91f.� S�[x�s�a����k�e��|]�'a������"�U]��������˼.�������R8��Ƚ�KuM�����V�Sˑ3��a6nԄHY�:b�Q��c�Ǻʁ��B)�I�5b�Tw��SW̑�.}VƗ����n�o�+�4��&�\���氾�Zv�^�T��L�0��,;\��;}T�6�'J��/���`&�[��{t��F31V�����J
6b�Ȍ���p��zm`�n�:��X~G�S�	��@	B�'L���"�0\:�Z��4��4RvӢ^��D=���L�҅�X>ܰ�H��.�k�v)YOI7��2:�ɄJ0�� s_��ůhu��r%�'5��N0j�(�g�Kgݤ�l@Z�M��a��u�V��hF��J�-�X��9d2W�l^�Gb��up��RVs7Ŵ���D�/�D�D��zKYMM���gi,78���؄)�U\�jN��-89����$����W���	N�nM�0k�*'�or�.�U;f���ZN��1�f������а���c8������a�m}.��I�M&Fh����ʁ�.������Ѹsn�%��Ό�aSѴD6�愃#�M���lrs"�I";Jݪmfй�$��uk�y0B���e�,�91�Vs�K3f�lh�~��1k����s��-���&b]��{9�C�����i�f�]�Wz�_�icf1'9u�ޗ%N�˫j���p!�!�&Lu[��RZ�L��ԭ/��w��q#�L�/�-:�R���՚ߺm�2�ļo�[��0b]
Xo[t����	Oz7'ѦVlY��,W�y3���x�&�}�zR3PS��i7���C�B)&u�B���b�)$Rs��٘�&p�S�u�`��@�^���&f��Y�d�Ժ3���@4d�$Ѽ���f�Ǹ�.��=aWD5�I���Y����lAK`M��5�&p"�-�N�2�vK��Nͺ�y�!U�Ww��13�(�As4nvmc�Z��� c�&bYҢY>��������ɣpH���8��m��"N�@mJ*H�<a����� ��SZ�z�_s9jJ�Y�7�q�\�f�7s�"�np�6$�luN�8�.a;4c�olԄ�Ό����{��Us\/���9)����Q��(����(�� q�L��a��+�<�,�,w���M���^�K��ՈI�ui�X5���ͯ[}�Wz�����n�A3�nf��@�(�s���d���	2bV���:�;��`.�8��fpOFNĺ��B�4��t1f^�Y���x֗Mq}q���jy���گ�SU[����:LǰzI>��s�V�`0��Y41H^�nNU1�4`�u�Wsx$3I���5	�-��/˃�R3v%e?���3p�Ѵ���Y�۰I�����*.�e&Mḻ́q��yj8պ����� �[|2˩���[5{r�ewo�G҂���~d�<��I
)J�MQsP]��&�n�27�C8�v� �U9��غ�]7c�VRι�Te��X��U9ϧK'��51Сf�Z��P� 0#��X��h��|V��F�luHZf��N,�U\I1'8]�D�g%/�8�7O��cf�^��"Pہ�
�/O�dQ�1}��f�s%Fm8k*GMi:�7r��,��]{3586Wd}��b?��]Ϋw�%������[P�@�KΡ�Z��9I�N_4�������ߨ��f�%A�����x_ a�κ!m2}�:2���`�15IH�R�>d�Ͳ\:p���{��2w{+
ƌ�$����kASs�+������e����Ȅ��bY�!s����3�8���M`Fp�(�Zp�l����t¯(e�jU���˦��S��[WzU�)�qYLl�)	'�F憂Y�G�J��wI�Ժ��RQ�fAZ4n��	�����Yi8g���[/4C2`*�f��,4'��_��
"w��]����m����&6��r���wG��!*.����/ĭ6��uQs�O�H̵Y���4���ylVL��UTsoͰA����rh��k$'��{������Lĺ��U�sx����������#S��U<.�� ,	�kz6�̎��ʮΡG΁,<u+kf�_�v����^�Y���)�pa`S鷲g��ybҲW��Ͽ$�����-�dV�L�F�[p�䨑�&�ך,m6��p+�µ5p��Z�����T?�\
5�2���s3�Ն��	S�+� ]��wC������A>��Q�N�ݺ%I��T��Zd��u�I�f�sn�Y|d�N��˸�uBs2��
`���&G���uYhg�ru�n�\Mx�Gⷘ���Ss,�IV�.��F�e�����5i��(e�������İzi��1K~�U�YE2��uX��c�Af����T�"�%X����������m�<Gq�.�/�8V�׹�s�����Y�$�D�;��\�uZ�q�^X�-����:u�54����1���Ȇ�r���D�K�Z�FςC����16wo���F7�N'D��%�_�0�b�m}��4+y��%�dj�uY��|�^ףu-|ysY.K��u�\b-h�\��V�����28d�U��<`�&\u�C9�:���[s3S'�)[�Ϯf��i�.[�b�\[2��M�nU܀Y�`�9S�d뵏��l�$|;�'0�3n��2�Q�X76��H�|��4f�nM���٦c��R��U�ufE��뵴d�%�f��A9b���"s�sIb����Ԫ���&b]��ͱ��o��^��+���$3pN�����̀}&P׹��9=��+x� ���2lbX���r�lxEj�&ج�f�,�qt[rV�0�������o`���U_xo۱=u�?rլ��\�rbܗ����i�Wl�a�=��}����F������:���62aJ�A��~$4��M�K0GBҪ���m���ubF��-D�V���e�$�����Huw��}!ƨ�����\j��%z��'Sg�½����S�Bvc���!N��Ӣ�slmL�뾖��~\A벍1�����V�Y8,I���OaN����'�q���`f�YDd�D/S�	��@	B�'L��,O1}���]7g�rG����ڴ��Z�j�b�o3@���j�|�S��_�fj��Q3���RPS�6�˃�r"3`!��D�{���؅M�����g���VE98!���l�< �%ƌ�����y���1'�bVIΡ�X�G['&,u�8A��xk��]t�E�/̂#&h�Q���%1a��F�<�c�1*u�'�Ѵ�ud䬧�u^�׺���Z�<�mɈ�� *2��pܔ�A�M��̢5cf�,51ul���f��q�.���� fE��!3aJ��̸A�D��+�u��̢_,Lu��]�ȌI�"�Eg�8KX�Z�	��m���ͥIz��%�f�و�#�M�u疚����u��S�̷d�ɍf]O)9��RV��:�Y>+�&bYIm��S���Y�����Y:k>����[xԀY	3bb_]�(
3�����}��ܴ5S�kf��uj.�$̊Yh�9��,�`̄�n�m�]��&X��=���b�Lf�o�6��������*g�/��2��t��Ь���I�M8b��W�-Z]N���F7|��)�-���pW�1�1`�$a���ڽka��ݓ=3j6������l	��Zv�΃�A�����4[�)�ǣ��}O�uvo��l�b5�2X2p.�31V�Y��j�͐Q#����f�Y�`԰��[Ή������RV�?�q�H1���󩻁G�p$g��Mr�i�����eg��d��6�࿷���nYlu��,�uJ��N�@�Mc3�%�/)8/c�$�G����aTML�A�^��cĺ���Yf�|�A��`���ݰ��pJ��.��Or�$�"��Bm�$[3��0��'"�3jp�-���f�HRs�U���2'�?Ʋp���Y-fq.����l؈��[9b��g�4�Ű�~0���8�Y���	���u)�� �[�l��)��k�4>���|_�O�;~zŤ_ �q���L�n��\8frsj5���~DVI'D��%�_�0�r���53@����
e3Q�iSG֨��"��f&�.�!�岔0`�Tw����:p��Q��;�߬)��s<��3�Irw�٬�'g�fwl�D�9I2k�8�\9p*9W���CBRT0vI�VWO74`䘹�r�������<��^���fR�$��p8�ʨy�+�x��]5+��QaL){R4p�,�u�C&L�O65���)�
���9�����-�ϸ��Ѫ���"��B���T��A6ܭ�\Vh��NL�E<hp#F������Ĩ��)LF�[jd~��3bb��PG�ͩw;�|5)�"�]p��ڲI�;ul.�:/8���f�J����Š�)[ �́����Ԋlv�6��ĸ~pds(8R���Q�R�O�ʂq��Ǎ�ev'�ȉ�O�&s��^l��[��>b^W7P�f�l��_ ���q6n�$};)���ҍ���͙<��!C���r>+/�b��]�`��fuN��=1.S�y4Ϣ�v����:����r�D��д����1�H���w���<8�Ճ�sE�����%_�[�ͤ�X���̺���R�u��s++�N-8f��f�v��5fVo���p���f�=���zݲ<uV�l吘A���zké�p����j*�\���v3nb�g��R�W͊�y9��r����2����ڞL-[[3��Q~f'|�P�f��K�<���h\�����e'Ÿ��j̤|�n�R�k'b]J�����3�ᬋ���US����{��Ȼ^Г�Y&%�
:ĝu�U4+u֛�W�Y}9q83�|����*\�3� �4zU7-gٯ#9�n��R/����+���-b4g�:�]'g!��$��cٓ��jN���ߥ��e���J�9f6�fq��ˎ'7���'��Q��Y�w{ݠ��ck�loF�y�����zj�Y�h"֥Ⱦ(b��#�)���ͦ�`*'��̑�&LH��Y�\+��0���f�̕ܮC'D��%�_�0����P�����͊��,XK�Lm�Ԣv3|�~�W��z�F���rUy��½`m�>�IhgM��D��T��5�}	���=�Qt��gS�{���9iЦ�|�e�Psؙ����w��21u�f��ḉX�}[��b��1F&L�/ݺ���T�v���z,�5X|IB���as��eg�ì4I��V�R����u��j��ٚ�\j������^U;y~9h$�G2�6+�&�I�،5�cfWMM��wu�p��fb\_�Յ#g[2Gq%��-�uSs�w�L��n!Vs�U*�:2_4��d�(���Y4&O57b�ύf��Hu�A2��/��Q��Mκ�'��'��'�r]�h��.{��s{7"Y���K��]�p�9���X�6�z����PY�+��Mxһٞ��]8�}2�a	-u5Ia��dΕ�S��,^�{�4cSv�ù�(n/�-̜�� x��r�=2էv������,�6�[�=s_�z+G�E�ȗ��*�y�Rrfb8�|�y�FL���;_�f��9���ۚLĲ���Q�d���S895��s��D�e��8_�u���(uG�:����&��Q�ˊͽR�&&��꒹�l
�ؘ4�0db�Z�uXX��f1�d�!��9��`N�
���H&&��Hf�f�M��]5��,k���e!掓YF�����$��"I�>��+{6��kq�Z��c`:J�*,�e�R�H2>J��������K��	������[,�W���r^$���ʿ����뼼Ьh&7q���F��|��ѷ��P���D���@m�	sW嬎��	E���� T�~y�$k���>�p�_૽�Ѭ�[�6%f�V��szY-Z fjh6l�c́@M��kc����J��é�΂��&��%&Y��:�κ�Y�*`������m�M��j�,��^o4j�b�� �2n�$һ��3�2f
>_�����&)�s��1r�����ڹ��L2����M��� �+�&�~Q-ln~5�.�u���$��Ƿ��7a�#�|��u[!�u5d�]�����.�J�!FM'_���R?��^N���l��!2�[�es�O�ϸhe��%&�u���yLo�~��M]���@4lV����[��Ȏ��A���\��lq�!��	��Ev��9䉩`��p��ʵ��:9b�Hպ��s̯����I��n�xZ~O+�N���u�]����p��p��ʉ��ͺ�9��EP	Bf<\n�lNL���V3��Dq=RY����X4`(4��1sl��5�q?�|a8|���_�
g��9lݓ[&I�sj�$��8p�U����pĜ9�b�,����kS7
N�3M��f���º6	�]�d���c�;�Ȭ�j�i��:4�vH;SցMĺ�߭Y�O�����,�[{�](]��6�nW�Lx��k7K{Q.�W�/B��z�Q��I�Y��8�V5]�@�'��dJV�p6��}bUT_�d=b����[�@ز���u)�Wa!=�5�I��x��P��ʛ����ż�q�'��,�E�x�ES-:��|�gC&)��q�rWΪ�q�ec��!�O֙Y�+�����D�@���&�����h�p�.d�v�p���,�.���̅��m�4�?712/��M��k�mw������;���+b]��Q���ğ0�7�f��`Sr�#��]n4w(Luf���]�r�����Y����I
����3����u[��B31>8��@7&jY���C1�<4aJ�~��{�f�ֺ�0sґ9Jc��V��}'xI9K��~}���pи�s*�������G��h6qW�ȑsYԔ�r�\�tX�u�8!�(A� ��I����>�p��稛��ҁ��jӦ.�s�Y��Z��K�6�^GR'sb/2��$��ɦጣ����P�[ZE�'�ݖs������ą��z�$	u�̀!�&3z٢9��ԨIr]�5�ѷ���e�707|9����$��p�df7ղs�p��jbX�^����Yi5=э^����f��V.��1s���'�z�9��var}cd��R\!l̄��ͻ9���1b~��đ��[�Pr),PfФ@��9f@�����qA9��!R�,ܸY����%I�(u�,��ߌ0bb8��礚��.�s^_�uA#FM2�"^�4��ԹY�eY�92b�>tr��g�2�R��Y�M�5aJ��e+��Ͱ����y2�[��;Z��[��������-B]ta�3[�#V���[�/$��n�L��Q��<�1s �J0k.g]��VN�A���a��$Y��b27"�P]9�f	� OO51����j���&<B�Ç�	�1���A�0�rj������\P`���/Ԗ��Nх�v�)#��d��4j���R~�9��pTD�S�	��@	B�'L���Y.b� ���[�5<f����4p�f���K����,@�.hx9����/2ˈ���uM���3ڌ4c�3�H��Yo4K�Lb#&Yfj^������qs�3CfC�"�F�m.-�k�r{٢y�u=>Sn�n}7�fa�s]���ਙ�+�x�4EO�2����F��>��w~�k��)#s�����Ѡ	��p5��B����Wf3���"��fO��u�&<���s?�l�Ԅ��������aJԜ��L�����F7�:n�Tw�`��v��/B]Td�N��k@fw��	\E�[�0_I�G��b��F�SFL�s#���LN��u=K��E�&�90d��{h4q׭����5�u5Cu0r������G���O݇\TW�L�ғy�����'g]�ufs���Rw���
^޷N���o��q�\�,��	�����@��Ct����<�R3F�4lb���U9�9�sl�������Sge�Thz��C��SM2�A��9܄�C�p0��4�␜3z��vj�֕�r�2+y"�1�9t��,,���9��a�,�$g��E��%]���:�rqBj;P�PA��	�, �g1}���­�"���U�3 V�65@�̷]��3585d��w���W��q6ຮI�9&v�\hظ	S�ʭ�Fsd2�\�N�L�n#+����B&L�3��
��a�[���,���e��b�@,M0jb�/��sܑ��&<|;-�f�l�S]�^�d����c�D��"��6h����� 1%���_�C���&�G������嵜n�Zm_�{p�籙�kQ�۾,̠9���͆À��uw�����.�1��Åi�X�m�t�5�[�L�Wm3�F&�����0��STN��Y�e�0��p��ZȞ=�_��?��J�I2|�e� }4��0��%�l�,�8��ɹ�%�RgB��*-�au�u��u��<V~Ţ�?80�2f`Ą!xԺ�,;�7{W_�0Au���'��#nw�W������z{y��Fﮉ��jЄ��Q�"3vY�9h�!s�	c
5��0Nx�>���sE�'�1��Zk�̢��7},-�7�&�Z4W�͋̄H�0G�6�6IF)3s�9�?9	mׄ��[�jĴ�'(2#�X��[��r�y+��,�[����(�07p�tp�'���=f�,���A�\z\6�|[91�]�庐-��C��ѢY�Sh���[t벞+v̅�#��.
c̀	9ƚ�r�oڲ��FN�\#�%�O5j�`뾱u#Ѡi��,9f���f����9PozK2r*y�l��{f�ul����BU�}UO�E�r6)�^���Y�6u�Vj�yV6`�!�L��� �u+d٬�Rwc�L�Q�^u�n���N��N���	��&���������έ�X�"�L��Y��y���uٷ��as��j��_�W-a2gpq}A��̭"�&�Ό�;pBH�b�nvc붐��a�Y� /�m�Uי��#��C��_o8n��LU�L������H��f�,��v(j�W�eFf�ٍ��L�Rd�hl�Yx��aҽ���lm��D���O�e�̗G�0�s/���wX)��M�#�MɎ������a���������"խ�*,�d�˯�������	g���E۸���p�n�e��+�P��o�,\�~�WH_��u_>��A�M|�]Z�
�C��}ۋ#��HVc{9M?2��Lj��Sw[^���+���-\\���of9߉f��D�S�	��@	B�'L��,������Bs�f\Q�f��ڴ�#n������g�?cW�!u�)_35)��c_M/��gy�&7j�?&���D�Md��ۧ�%��Zw�-.2+p}�$}[�������W�_Wͱ�LRp��(�����hjݲ�s�] ɺ58���%��u��e�L7����1��K��ނJF̻�l�>�l�1r����<]ƫ<��I�"��9���� �d�O���F��3��:�_k���{)�́��J3�w��0j�dUcfy*����8(�]8�U���$�����`&��j���� �&�uj^%�ָa�Xt��5x�d�����
�l�lv���AlL�*���e4�U�S�d_Flb	�
�0Ԁ��mZ�M�Y`��I�a�����-�d`<EF��c��Rsalt	7	Ȭ߮���:60&�5p�2C�&b]���"桖��X�=�z.|+�`�5�3����>{��̜p�'�(�A@�:0l��53^�@����N98��W�ufb���a3Hb#&b]
�fn���p̆)�B�R8AϥZ�'��":o�+J��պ�ny��B�FM�˫�>+����_��h�#����ʁ9�ˑ㦤��_�BN�O'D��%�_�0�r��.��u3�]:�eMk�I����r�Y6fj�E��z�uZ58�Ks�t&�y�}����*uKk��K/N��z�������РYjr�5I(5�q�7�\��-[4�ƌ���$��܊��G��uٿ�p_.pܠ	S��͍8����-���uVêus�]tb�!&���%sp]w9ղÉ8f���"�~�#��C�I"�Mx\��z����j�	���}��})�	S��;闢���Z7��G��Hu'�9ffb�8J���`�,�pfIֱQs%��r�&D�V�
?�Np2n��Rw�>�,~3�f�s�����C8�Ju8�z�n�`�&�~���Aky�}׹Y�mY��H1�/(0�f�54�r���Y�f�=	Ʉ)�ʮ��_��,<3���FL�#ԑY�M���+����E����t\�q"u���X�?��N���`�&��xg���n�4��$Y��n��1s��!S�:0�5CW5���~�\��uy�	����C�#-�ґ9�t7f��9	������S��)\����6��.<ed�^�7�ۧ&ɡ(u��̆��5�����C�8!�(A� ��I�Y�}��P.��Lf���ڴ�j5+���f&8���掁!s�M8\[w8��9���0������#�-�jf��m�k]݌`��j:������;��uK`��I� ���+�|^��M·��E��Y�
�l�E�٬�����
0hج�8-�u٬̢Zfb��R��U�u��$��R'�	����h&����r�pr�m|c-1u�s��́&bY�m#��_�Q�rr5CN7r�6d��V8dnUr�n�Z6f�E��8l\�˛L
"�j1pЬ�z�AS��2��+�D��߫s��l��5No�����9��'�c���G���ѸI�u\_'6�s�W�_��aν���f���ƌ��u�}0Kҍ��-e��7�Ss�/��>����cH��[�C�8]'f����0���"խ�*�ټ�kC&�~�����>�P��=�z����-�:9h��U<����8S�bV��J.�d���A���Yp+�l̬�AM\K�����>���,��@2s-�պ/*2����V�[1��Yw0K��:�A�N'D��%�_�0�������#v-����Z��C�6mj�Vb�n+f$b����r��S|<%�t,�3H���0,2�\~G��L�-��~�8tBB�n��͡�,I�"��.�rpBP����y��s�����+5Ku����\���x�C�p�f/i^���ub�RG�0��E��d��_��.�a�ڇ� �,�M�Y3f��b���acf`�\!nB�n@s��9�%�ܠ\.33p�4ɷ\�E��1r@��Ռ��p�[�YLrF��:4`��Yp�,[��X��[A�뚢qsW~��S�,g�MM����.LjZ���m��bZ
dF7I��Eg��7��:�V *b�Bu_�1��R$9B��{�;��$-"�f#�k8�y׹Y�Qj��M�-23�gk��L��������Rvc��Ó���fNG8��W�9ݐ)�Sw��-<�i%̈�!d|]tY� "̐�6!	`̰y�07[M����R�fԨQ'	�bȍ�wm�n��6��l��X2M�-%8`�,��'E_w3pBﯜ6l�՜�w�L�l�i���?8��X2+�fQ�� ɷm➮��d"֕�`��9O�FΖ�I�>Kk��7�J�#�&�1C�Dz8�s�/Dh�T��l��T͕O��3H9|m�M�����̃�A;'6�xZ�W�V��];'ɲ�eݷ�fl�:9+�����X�F�F�8����Z�5S�90j�����[�pЬ���u������Z��0�Ws��,���
'���& S��ԐAg��J��qQ�63qԍR�,��f/�uJ���g���=<&�-��,��;�n#h�&��ԁY�qZ���.�ϑ��r��8�IFͤs�ɸi�-7`��Ǐ3ɺ`#f0fNi7a�;��ӥz�b�_+0���V	f��j5f�к�����i��Y��S�@"&N�j.�%#�
mi�9�9D.lq`�lW�7èhu	@9��1sMŐ	S�e�,֕<�U��g�鉆ML�ew�ΛubS�����(7Ӑ���g`�`����"Pہ�
�/O�d9����˚���b�W(��:M�:Ҏ�mR+�̄��=�uy j�+K�����,GM�/2�wK�!p��Qp�7'������ֵuSD�������	����-���+�=�����y��tٮ��h
7�lqX2s�夐��Z�efA<a*�43��&6��v�EsB�!8x����r����@��6���9�q�M�ҟ�W�9��s~�9�I��82��vŪ�oW�&.P8	��u�ς�����[�uZ(Ԝppb�of�n֍�3���_�QoS��X�t����$��R�N�xd�I��n=V�/g�"s��f3d�59��MZ�z2ۋASu��u�LS��Q��,��'�����,�U��:7b�S۩��Y�[?�p#'韜A거���-��s]ļ:���}����3[��6!&����j�����F���������Z�uz��B�l=5������H�p����d��&���&I'9����?���u9������p�?�nt�����d�Ń�5?��	Sݭ��]$fR4G�C���A��9)�_w Yo�9��j�N�B�xؤ�}����p`vٖr�j7����!�怱����Sb����:�c��8�Y]w�lr�m�Mzj�%�dh
�,���]tGN�n���Ӭ#5���f���1T�Pw��y��u�Ĥ?�_C4��L�;���uWc&����4�j���1�.5~����t>�Ą)�F�6�f�U��[��#�FĜ�g�
׷�lx64$���z����L����LԈsV=w��\�5Z�j����mWo����^m��*��q���X�iy4���@�N]l8�w��Tz-{2wS�I��R�حB�nb��j� �5D�Nb��%�P��7���'�ϑ�>ù��M�#X���-g��"C�E ��9nVMNĺ�Nb���=L���&L�Gh�9�CT��c� �l 2+�$Q�ާm���x3�ęm�O'D��%�_�0�r?����xw�?,�Y�pV{֦M-27���ѐYi fj�3��:�9�nZ����d�z�5	�|07a���U�屩�y����;j��7������S���Ig)?؂	F��4e�z.2���!Qw�<����F�D�+��YK�/#8j����qIr�Acf��1���ۦ��]���?��]4IȉV��cb����U����KM\��'F����r��!9IH�d87g�t�O��5bs�rJ�U�����7�tMξ�uj\ؕ@���Z����dz4p�ka���t�x�����$�ʺ��f9Mݩ��(��lb���0Kf��:&��n����lp�,_�x	,�u����,���R���6�|��R5�²&�a6�:0�麂���D�K�^��=2�b������ʒ�Kh�j�Bss�P����2�25��N��S&fA��fV����L6s>ǁ����͂x�tS}Z��I堉+�!���ss �e����`b�s#V��Zxmuy��lD�`�L�,R3b��˥"f���Ǻ?���E��P��/�e��xl�Y ��7�I}�����Y��+�f�i1p�΍�-W����1p�nS7��R_{51����r��TS��h[���L�e�/gc+�f�Ժ[���pb�tC킻Rh��r������y2�7d̘9�pJ�!�J�9�$!��
dsR�o���Gs�9ђUfܰQs_mj��p��r��G���7q��)�Q���B��|�dR��;��Y���V��ai!Y��y�,���9�/'7�n]�l�qW,���i�^�cMĺ����Rs8�S!+�ِ9ԩQ�8G����94r
GqBj;P�PA��	��M/1}����8l�KfV�rX��ԦM�Y���̶k��� 1SC�As�Zr�����\f�CҶ���/��N�NW8��q��I��?��M�)�G΅���=�$E��5|���؉g��!3@�&����:-�l*Ϸz��+� �IJ~������J�e�<М�bܘI�9+�"�!�R���P�j��7����;F������C�Dz6C+5gȡ�L������+��qA��̬�������F�L3Ǹ�6���k�:�.b�����N�N/f��G�������"OLo=O�FL�}zB��k[��U���L��m�P�Y(�$�Tg��М�I����}Q�XM�ˌ��X��2Y�LW~�J���f�K�&�_��m`�<���!Y���i��̦ͩ��q/�2��Ɔ���#���bsk�٬$���p�On1a�q$�#�Ea��z>�9-7���\j�$�'s3���΂�sػ'j����٩Kf>�=d�U�f�z�������΢��k��;k�p���v�-�r�wmG�MB`f̘sZ�7P�G�l����.ʦY�#�f|QӠ�.�w��Y�䬌0n~��Y�Ka�P�M3@�Ž��,1ãpԝ�+p�6�Y6I�G�C#g�\1��$���Q#���v{]�lg��IN��lry�9�k�Id�@��&N��栴�CWĺ�chԀ��k&jYN��v����SP��Ǻ�9�I�D����w]��Pssؘ�gI�Ѭ��fu��m�؜-����CL�1����p����u�&����5�s@�ow��GN}��0���N���[���ٸ�1ͦЌ�N�氼+��51BZ�MK�� %Z]����s#&\ɯ�B�hϋ��ܝ��)!Q�6���Y�AL��Q���uS#'),3���<YAȺ-�U|���i�F�.�kO�[��)�2lN��FS��܃峆k-c��,{6e6��4�ԃ�$���h���eS�;�9������DD�x΄�\�S@���)�)��v�����&Y@�b� ��>��n���g�M�nΑS���L����"Z�f�T������$8��w�3�FM��-��~�҉��-���0_eY��D3�w�$d#g����`
K�ͦ�Ė.Y��.֝MԺ���-���	�&L�7��V� &GLq���F�İⶨ9�v�yEGt�O�'8[���WF3����L��_���&'L�?+w[����pY�d~lh��k�H��U_��<�[�eC���4)F+;��}0nc)�E*���b�̒Ti�ׁ��{�P�[�n6ef�x���Rw�����5����Y����lV�bκ�ur6���g3�=�¦nM�,t��A?�χ��)k�Mĺ�N`����j~Y�^Kx��}��!s�ݺ����6�97��#�����/B]�wE�L���q.Bݦ_H�7��T'��F̀Y�а��?�۱8��!�p��5Qsx�a��?�[�!�L嘛�������d�u�sP\��j�#��:&�YQ0l䄉c�.�\.\0Q�r�M�]�f����9�3�bh�S��U^~ÝE��T����>��,�I�ŋ^��"Pہ�
�/O�d1�����0�p�q���,c8P�iS��hە;�ײ �j�>�N�6�݀ﺦ\^��������څJ�����]zK]L�΍����~[�]gf�h�,��e&e��~���n�>T�Ƞٌ�uEs�M֡Y]5p6� �.�w��&������W�Uh�`*��v����s�)R��Iq��L9=��}=�efK�\</�ݬ�EY�'&1�q}}���P%jU��X\~+� �@aJM�`x`Y�u�|V3\�~܄��$��`܌I�"�EE��ܜ�G�k�N��mz��xq$	��ga]�fԀ���3/�_��Rκ�,#1j���r92d�M�mj��Y0h��IN��
'�f#'b]J����Y8�I܈�¹#Yxf6��ln]��Q�Ȭ�:-���%�.����@9h�80��[�/\���:1O�D��+]j�,�Er�-�R��h�À�$��u�ω��ꪩ[���f�&�|���hV�ƇIhl�p��������(j��PNT���'�z�i�DS8�f+3��a)#sW�o���T�����s���ڽN8��"Pہ�
�/O�d9���c���Y����gZ��e �6mj�|�n+f`����9�!W�9�F�as8�k��+y���[���0թ�&9��Y���bNW0�~�Ό�%�̛؈q��h^p�wש�st��<�4n�0Mk��W�3��d���3�����sP�N�1a��`8�|�[Fp.�d݅�f+�f+9�I�^X���$�&L�����Zj*ߣ�ZbB�Z�y�YpWP�{���k��fnE(�n�Q3p��kk&D��7wwAY^I���p��^5]�f�[�L�KՃ��5���W���s}�k�`������ƍ�1��Nx6w�!�Yҿ(ud�����8f�^bl����f5n��\Z���-N�gfi_�7Lu��N4�M��XP��o&|^��.�+u����(u�Y&f���K熉!"u��&KM����Mx�����n����0��.2��]j���Hu�����wy�y���0\�YpW��VMx�T���s��0�?80|�d^����\|�kN�Nn�&$s�V�q6�FM�ԙs�W��|[H��Tg��sV-u2r�/�tkv�-�����e�L֭�ީ�p�q�0e�BglǆLף����fw,$�N$1�d�\��sO�%_����u_ǣ���E��k#�d�$غ?�z�Q���g�܏T��f���7�e=�9�9����#��\��	C�ӿ�,�B8���9Z�����̍�{t���Fҁ@��}c{r�$뎸���*(��J�9�6�Y5ud�7���Z�j�,/6`�!�L��{`�p�UbN��Y4f�E�Q�^u�n�f!U��/J�mi�9��4\��w��`s�Ŵj���Ff!�$qu�|��Z9�f��J�wĒ)=�3h�m�1��A�5sHM֍?�236ֺ��z1��md�İ�B8�r˪����*�#7h��F�xy�vS�;d,�x�������V�i�n��,ݛ�<Ѹ��>��}��Yw1m��]4ì{��; ��?�Ġ�X�rn��ܧ%�Ԅ'=7�N1�q8��Ă�(�Đ3��^]'f��%�[�&)�Hu�
K�̒��p?R��gs�G�I��ĺ�9��� 7]'g���*�{db�M�Ƕf�B>��wu.J�_bf�C��:3�����v?�ɬ��t#��j���*-�M�>V��54jE`*��-��"&��fY�9�.B3��qBj;P�PA��	�, K~y���#|���Z�jk��ԦM��Y�ۊ9�W��|�%}��p
��LMy��^��*8�.X>��6�9H�I��B�ͻ�h�T����9�O�ʀM��忻b��cf�ذ9�Ѡ��p����7s J
p��l/��)dX�dV�����$�}��7��@a��쟙��N�r~�Y�h����b�7�z-��$D�;�����^��/J�9��zl�K�'f`�^���*�1+��I����\�y㔍 Yj��1������O$GMĺ�c�64ǌ�� ��Ku!:���WSӿ�r3�}�%�ƽ��gT[v�.@aC&)7�e�f�.�l��rF3lc&���/�b���4[�n�~,�W	Ͳ��n���9��s�WWN����鵍�"���t�,6#��/��_�
�뷻|��U#44��r�D��������#&L�C�ceؘ��:�����Fs��TwA��:.F1q�G��FΦŜ�j�$�w�Ѡ9t��*���v�B31?��,�36�R�ڀ��ݑ#&L�'�	��9�I0����É�&9ɦ7�̗ �Zwڍ �ܮdr9�ԁ�CN��z-c4b�\pb�T��G�-%���VlN��FN�O'D��%�_�0�r��.��u3�]:�զ����#GȊ/����ـ�LnM?��,2��$8�9(�v4�7�R���{��o�l��]7�m��qS[ .L3d����Z4g�9r�F/�54c�@�\��>�76p��f�D������3Ι��hV	͂C�v��0}�8�m1�:���,�U�h�n�I2�ƺ/�j�����LxX�ǫ��&����_�]8�1͑y|�����$��!��ˆM峚�����h�@��$9���9L&�4J���}��Y��$�_>�}����S	u�6f���#I�(u�Y8�ss�#&�SK������Rκ����Mj���tac�n�y-���^�5��L�'�&���h�D�K���r9A/��0�w�c���y�C��K�?J��[���6����/B]t��݌�g��0�?Jݲ~!��r#db��R��UXjf�`�$���f��r�v2�r3jجa���f!^8o�QQ9��u���WM2�!�1�b2��z��e����	�-��i��D����E6�1l2�Ni3��wX��?97���I�"�E�7���-Q3N)��v�����&Y@���>�ps�-77�df�� �M� Ws�\�}陙�p���%-f��f`7������B�{�_o3k�ɬP9f���f�^v��9P.)7��I����!#'�����d��C�����@��pм����_[�q�3��S��0n~Ѩa�v%ӳY�G���Ɍ=i�0f��L�Q�^5r"j��E��뵀�G3��w=6,� ��έK�f�%�����iK#�e����6��&<�o���pRf���>�ܲ�L݁�4lN�Zg���4�a�z,W4�{�+�^66����d�f��b��T����l��$����-8��Oݪo�9��8�qsdF�u'��/�=8h�Y�"F~4fnŒ�~l"�e���Y�Eaf9���C�U=_O4f���y! #�M��|p��S>��C�R���^��JF�_Iw#��U6�s��Te���R_��[�ur�4��Z�+S��j�`�����·~1h��2;͗#3����f��Y�m�c�t�,�p�捫i��Y�[��͉a&	���O�I��׭[�1F?�#�1j��)��v�����&Y@���>�psĭŢX�����C�6m��<go��k��za�3�{ڟ�qk�&����~�1��(g�M�1f�<$7�������F��[���g�DY���EQ
N*������ܘ����w5�bQ��] �9C���4/J��:1a�#sU���2��/�u�ſ0�� �C�R&�nr�q���j�A�D�P�P[��nD�:2����5b�G��[�mɈ�� ��lM��~���3�1#��I��%��?��#�Lĺ��r_�6xE�'9aJ����/ 55����-jZ���m��·h�\��Q�3zu�h�ϣm�ԑ�Ylz3h.I���] �X7G���ud�b�w�Z�fs����6Y��V���ऎV��̦ЀY�r���X�S/4�r������e��l��H��jO̝]��6�.��QfH1c&� ���ņ�b{Ӷh*wͬ�6k�F�8I]���0�mWN��Ơe�~˭�����%������zm�fY��`Ff�̬� '6#�5?*cɬ����f3�
'�70+��6��r��X�ӣ��f�]�b�s�R���s�^[��Ib��$L^[4nn�E�Mm�̠_N���7zB��,=1�iP����Ԩ9qV�MI�<K��?\$�����S	 � L��^�1�\�����a����o�#��M���ux]��,���g�Y�m�'�0S	�����^s5���-j��bF�JE3`�{�+������j��S��(u��P�Y�=|��W��xԀ9|w�J,�f��0�&�n垶�&j]J2�i��[aJ�,��ad#�lq\64ϴ���e��]���$�1shS�q�n����uK�}�YX/��13$��qh[?7���F�4k7���h�_�bb����,��Ӭ]�j���?H���5�s|��7�@,g��.��0�ߔ�C����6k��M�9}b�ot���^_�ۊ��n�!/M}�7�p �*�8!�(A� ��I��^L`ξ���~��6q�6ud-�Ɋ�3�{[?��9T��n,�r�l�5I�9��c́����H`F���e�РA�N�Q���&�����lz!�Kj��J�sP��P����C�ȑ��b
O}4d��I��u�q��X�j���}T��}��嵮f�ϯ�@V����j��\8�ѥȆ��_�U��9��|�ur��9�6u!'�&����B�Ժ��2��̀q�?4G����Y`*��`sh���Ƥ_�峞bVL���Wb�\��"֝v?��11�G�#s0C�l5IzE�[�Uz� O�̩Cs(\�����6��C�41e/���׍�����z,��'��C�z�!3j�	W��Sz�[���@��y���42lFY0տ%	�`u��]\�*�;jn��&���f¨9�b��P��:�#�&��\W�L����5�|�\h�;�s�Y�t���Y��6�����FM�NK��M��0�~ĺ�|������&L��\��dџ�h
�[l6���	S��^��6�.��HuK��y�y6��D�Փ��#ty�i�Ɍj���&	+�tٽNf�T�9ޖ��L4pb g����_M6�Cb�k��,Nrjٳ�ԲWsn���v�s�͸���uߤ�k�zf
�,-5rv�em&Ygy,�����u`�,,k��W7����(��,GQL��l�� 2��W�]��$��uAsSOb5h"֥�ˑ3�Y'6��� 6mf0�Gq���?o�ȉ��ʋY�u�x5�
Y�N��x�6{����R����
�Yff.b��չ�E9j��n�ӣ�֩Y�M�Y11����[٘)��뽮du1��p|`gSRo���\�-b��LUs��Y`j��%�抬�5q�#Ա9oד�!N�#�-��[��hb�����+�L��g��yI�9D,K�s�����Mx�/V7���S���q=�؄1K�,\x��6\ug�3+�"��)��v�����&Y@и2� �����s�=7�6mj����)���|V�
[���j�4�r�<5	�W
�R�oZU����A\�zo�� s��)\>��<���An��C5�%�d�t��[�dIϜ����������o���x!�>aJ��o������w���,M8l��Yw0�X����}ӫ���He+���|�x��Qs�~��K|�ϩ�xU��Xxn�ⓓ��H�l��5<P&�(/G�XRh*���`5V"�u7,PMu�̡q�A��&�~���ɀ9�V��kv�/T9I4���`��p�4=N7bଠ��&yʎO2t�-��(e�ʹ'p��cX(��&�Q�r]�6����p,|{�&A��uޠ�����ȾC1�QCf�e�//3Q��]fh؀��pȄ)�e��h�f�T��\�%Df�'�sXF��p9�������4�)[���ֲ)n߻�<?cAf}���ݓ�L-[zjn�=�+{��޷u�֜�/��`���97ff5��ܛ��፜�ߦ٨�e`�]��#i�q.�L?yذ�V����Et�s�~�ċn=.���R��,��t��!n��-�ŵr'֭���u��F���Ť_����Z�rf=���Vn�nɪ�qS�n�f���E�3����jٱ9��1�Wu��V���J��kf	�9��$!�D8�-�ln���xn�$az��!��xs�����NLLG�{܅S�f��ۑ�qv�D#7�u���~c�m3���j��a��o����i��L�s͊���S-{5W�S�.��`�F΢�9�I��Ϡo�lش�Ȝpw� !�pH'D��%�_�0����R0\�������Y��D#S�N��:)���Șb��F3:�9��A���Z�w�nbi7k�D�[��d�$_u�� ~�!
E�� {��I?��w��nj��>~7`b0���I��_2��B�z�Lk&�����^��긮�4�܉����Q�V����8t��{!6Wj5�T���V��p�'1~�t���qs��ɀ�$���=^7��r�D�g�E2�̂q�/�	���pwɯ��[���ƍ�p�݀u=/�m;��cf���@ժ��&U/��>�]��'�M����v��!s�F��z�y9�$������'�4ܣ��w0ېI�G�^�00�
�J��+ge�,3fb��R��U����N��n#7����f������YB�U�u��/IL�0�/�l�ȉX���｛�)���~]6A�R\1��ጹed��ԹY��:�)�&�<!�&��h������Բ��f։͒��ב|�.�����&bRk<�c���2�s�,�6|�?�Y�x��p]��+��嘉G��7y�.�E&Mt��\�u��&*$��b�5h���>�eA_^lbHFF��C��,�N����o)���"խ�*�ů�����>��<B�Qo_�-�s�q�uk�lV�@u��A��o~����
�`F�59�Ǡ]�3���$����[�%�8��`�_�WRLsnEWiY.��Ǌ�3��9��������l=����
����o�^��"Pہ�
�/O�d1�Rb� ��}��Ų�VU��t��f����������ڍ���M�_���<�&�,F�q�����������٥*&Y�f$?���I4�暂IRkynr^��:.��ӂ�&�*1`��V��uP���f��%Y�n�8d�Ц�lM�3st��Y�H^�e�z�b��E6|@�`�*�^��<vs�ν2�� ��9r�亙ucsa	f����3[�)��%Gz6\��Ư
2{��j��n��'���9'��r�d��ՙ9�����9K�}3�q�Ȑ	��s�fo$I�eK ���͉� �ph�^�u�(6��p�����nh�$��|>��lMI�fe�x�M����+pA0��n"������?m���'�������}/B2s"�_��hu�nn8bج$���E�UR��f��7�Q��^GfG&��eG��+up@�&��g^�`�.6p
g6q��Y��3f����'�q���ԡ��d���뼨7 &<B�̩���S?*_�f��L2'3QY�ӟ�w���LХ����O�u'��рY ѨIr"J]�*G�0f��	C�"N�@mJ*H�<a�d�[J}���xVsڬ��^v ��:�-�mW�
�e"6K����f��T>��,5n�� /��f�Y{9pB�N�Y���pb�u��K府�]g�ͺ����(e��Vza��j*��-9f̬+�q��8[�p6ÉXW��s��=C�i ���t���\:�㺦H|���4�r�c�AQ�:-��S}[��\�s�<H�?t����rȄ��5^�bV�n̈	����f%�,�7��������{��j�Pr^�͠q���� s��q��/B]T��(f�a��hu��Bjf�8���R��!�43�fC1�[����lp���Tκ��&&��/W3���b�9Znz]��P}�,X� #֥�[�?"�"�0�7�:7j�ٲ�6Of��ܺ$��ԑY�u�i'�&��E�����p�?Bݲ~�Ms�)Lu筘�o�H�X���a��ںq�97R/�&��k4���ugS9������L����,�0	m݆�_�b�ı�5s+�ܞ�1j]I/�>^�,E6)����fQ�A�]x��U��p�y5INE���o9l�27�bfy�G�S�	��@	B�'L������0�7n���An �6mj�\����f�g�f=�,���6|�uMr{=̼B��V�Lx��L�J,��ːtp�yɐIֱ�rl�'7aJ/�!e�ɬZ�����>͘�|Z@V �M��FM�ni�Y�'�J�	���8;��	LF1��=P-#8@R���_2d��/�k���)���A�FΩ5l�nt$��	A�l��ݹI���wo��`�L­e�m^���2�cf�����@��ey����4^�����Ss���un�4��;`lzA]���T�dA��y0�(Yw��-gu��n<�_���
F��q�$k�0�f��m ���r�,��]W1b��/�˾񶶅�f��,3h�,41u��RjNn9��,��t�ܸ�FG��βu��b��0Q-J]t��7k�2R�t��p2�i���6�a�1lfu���z5�ax���_��|8Y^c\x~���V�&<_�����2�������>�ɠY�CÀ��$��ա���ԄH��{y�`��3s~\�Žq9	��l	ȑs��Pmf-������:8�fe����8��:,��ؐ��z�.7p6=�;��/�Kq%Nf7r����I���ʉ�oٯ�r3��n�n����v2�I�u`��[`�'<p��HuQnL�1\��<n[�؄�50g��³.P����l��cS��>��6������Cs��b�j��%��:-��농��Ww̈́IY��������Nk�=����z��!�Lo�y� .��lj-�+�6,E7f������q��0��/J��'���D�UN��`نZ�3�|#�F�%��[#0�ҭ�{�lg`�D�a��G�h�f�ɠ)�/Kw��9��ԭ9�kkf�-�O�u��cX�L�����Z��lVi�:�8��>9f�W3j�z��M��!�~/��fجtJ�Y�g���t��77�L�joì{#�x.W5h三X�rn��v�o]9��`�,�Ǯ9�@Lq̣�Y�lbHw�ZC2������o�-E�^���p	�W��Huw��}�ƨw��H�ՄS�����J���,���,�� �
�3���abо
Y��z�*H��R9۶ݏ�����YV��#�~�p�>V�n����|�Sm=o��p]��-ɓp���$��u�8!�(A� ��I�%�<� s�]Xn�,V1A�֫H�6mj5���s��Y�|��s�T�^6p*��LM���8�O�1�w��Y��i�0I���+g�1�M���0rn�ʁ���Y��Ӧ����9y ��fZ�b������FB�n��2�=�B�ECF7�8$�N����L��u��{���|(fC&L���r��#��\ �u���ٜ��(u���?$.��L��n0n�.�dz4pN�	FM�-t�w�/Y�T�z.71�5�W�AmK555I��y�6�w�p'b]����N�	S�{���.9]���c�Aɺ#�`���G�m{L�D4l�$e^8ò�xuݴe��Q�D=<$�Vy�=��1Sd�Ig�2bK`5d.����m��|>0�%I�';��Q����u�̲_T1F/M0�s͸��k�v����
k���&���u�>��2���YFj~��9�tm+b���bh6q��Tg�t�����#Ձ9,.f�L[�9�/Hp.zA̺-�U|��$���b��r"֥�s�]��e�h~�N��9 ��S'g��ra�t������G,9bj0K�uZ�bH���#��j�a|-��dFL�O�W�v�)��9%䬅��"N�@mJ*H�<a��x�.��0��]:���jӦ.�s�As<�e�f)�A����w�qn��t&�Y͑>��Yg3!R�b���q�Lw`�x묦�u��Y�d�f�Z�u]ދ�4�E��3ftLry���p��j�D������T�T0d�ޟl��L�����Xg51�Y��x�݀��膯���wo��Z�s���:c�$ң9��u9'4�q}eVШ��[�	��h^����ʝ�aJ��{�κ�)tR3�A��Hu'�9��a4	�Q����D�0K��b<$��9�C�nY��f��'Kx�F���5`�$9wUؠ�|�,�Jm8�vV�Y����I.��B��m׾뎩eY� 1fbd�/fx7j��1�R��y�cL������{��T};^���J�;J��[�È��NA�k�Ĉ�bf�"���(u����?����N��.3`�c1Хf1�6WL�4���$Y��g�I9wS9��b�Q3�T�L�f�/�s�Z��S�Fh�l�a�Ժ�qsqV�� Mx��9��Ѕ��̱C��fy�	O�u'3 ��٤o��{ 3���ɨ	�*��v�����&Y@�z)����p�9h���Հ3 V�65@�f�G���Y�	��جˑy�_Hf���Fϐ�V3�#'\uO��8��v2[�13��6��26w��S��+4e'�X���3s$.��\� HWr�/g�&�ۂtj��aNe�ŨF��Sx���Cf�ﺰ
�W��Y0��b��R��U�u�Q��/J��'�9rd�%��R���<�sm�_�����M.x븲�'9��rv�%1f�M���,Hsh]ZdnY��n|a/�"���̃�Y�R��zl�lM�غ��U������Φ�ܒ�ENUm����~������x�x�r�V}���ɲq7)����ϻ�f��-�;gҽ���6s�Wo5"����9�aarS9=���f�kw���)�p9K�BC�ewMVk	v�z���3-I�E�[�U`�������Q��>��<BM����&G�禎�DѬ���1C&��ŅsRWH?eͬ��=��M�C�����5b�Z4fF��-8'ˣ�QӜ#�~�R�=~�����Ģ[�r�T@[�[���II��Fs�X��@2f��)��v�����&Y@���>�ps��"X�b-�6��ŷ�f�]�d�L����S���ޔ�$�6|3��.P΂��	,�!�I֭��y�Đ��!Rg��.�u�3K�.����('�[��Jf�_�D��̀�gZK8d�] �Jou8f��4-B��21�(#s���"YW2��+�u���0��P���-�!ߴ��c�a���33�*uZ+p�́&Y���8D�YH�4I�z]ǷG	 Y3�r�,^9GG��,f6r���ԑ�Æ͒�#gc`�D��������Q��b� �����gS�/�u[>k��E	Kݡr��a�|e��(u���jƧ�7lB�l��/�o_�$ F([h�on����E�h1.?4�7[@�oɪM��U^J�m���Ϲ�����"���n��J�5����_��H���^�@0+aFL��� �f�7c&��&��s;�n3G>�5ߘ8I[�M^���7�s�fe����=]�.����.y6l�b��Bt"/��i�Ȭ�����d��ZRW|X%GMM�2n�l̫�$�f}O����̘�ZW����9�g�0�? �>7�n5|a<��꒑���m��P��er6�g�&&Ay����f���-Tk2�ݜ� t��;Nj�*��s`�N���5^٣NM.示�����y|a�|%'����Es沉�y��]PWNM�.�w��F�K����]8�A��n���_��B&��^$j*a���I3qԍR�,��Ka��S��u��f���l�X��b��_�jV�L׭�b�R�aPM�����p�ά�u)���:�Y	8l��	S�eafS�3�n�\F4g�k&Y&���j��Z�Sv�˅�A5G����_>p�VUM���:$��q�<��^���/�uڱ�l"2p���\�fsSĬ�Jl�MX���x;�D�K ���]���ߤ�k�,�yTY簶�A�&&���9d�>7պUf3 א���
+��&�J�8!�(A� ��I�#EL`0g�7��h�����tK�9��=��3�9�~���s]Nug^�Ձ�y5I������/�g)���\/81�=��r��q�ƥ���e�P-����ԛ]���a����%�Jr�xÅ�f��Ҹ�rR(���\�u.�-`f�ĦW��#�b=Ą�_�ė�ʺI��;�ώ��@�	Oz8�}�p�,��_����f��&Y�p�+��2�S�vrFlVtS	�^�Y1�Ѫ���\A��՜�pbһY���h
�߿�QsS��X7fެ;#&i|�:2��C�|5)�"֝]���ڲI�;ufZV3�Xޚ��f�I����f2�M�Q� /��'�ϧ�)�5%q�6
�PC�M��rX�n�8�_7�8@Z���ux�����gsQ����Z�5:q݈����[��p�MM�F�齠�C&��� ���P̦��^jNE0�`�4�_1g�u}̮#s�W��FM�.r��"��ks�D����_6����h~ aA_���C��t�sqX8a�cs����-�fR�F�C�ʛ��q673&��#b�-pK��?u���pԜHI�F�17�æ��B�u?좁#�u9~�3�M唘A�՜�1C��C�u;�n]����&	r���2-бj~��s��>��@S���m1��s�c����f7��c�߂�9���u'ո��j̤|�5����l�D�K�_87榃��C���M���jW����8Z�rb�_���m���Q��1�Po]��B��1X;����3����*���.פ�kxl���7c�֝�k�f��Ĺ�FͲZ�끦xi-h��é��.��HM��
]�KlM��q��]����~�9��u�&&y��ͨq��ob�'��Ѱ��I��,s� ,�e��L��h��S���R:�i%�a8h�U`'+_!�X9Ql 2j�����p�Uwƛ1�2 3Ex�8!�(A� ��I4n�\?�p�`�f�\i5����M�:���w��J1S�_�]\6$��~il5O�FMB���-��1�n�݀Q��3�u�x�-2R��q�;\$r3�Z�C�Nuٚ/�c}#oL��qs؁3 S܎�+~������9�~UW�R�u��+p�ſ���$��\60���)�݄��̠IBJ���ZI2��Ô\��r�~��I��;���FM��g����IBN$�Xlܜ:�$ܸY#6Ozw����pw���h�䐘Sq)-�oU53��kBn���Nllyl�����9�����$�n�:���u$�Ɵj�W�g��Hu�Q2��1��Hu�v1�s!0'���uy.>4����'��x'��$�,�E���C����,���V�Y�F�!hC��bE�K�~�/��[Jr|#�qpr�S]'s��+5Ia]`��u��4ej�f�6�&�lXzP������<�@�ͺ<�]�W��m�I1C��26pVn��,�՟���J����r���%v6��ulج��7X0p�05���us����!��pE�D,ˌ_���a}�p?j�u��#{ۣ���Y����$&	g���:.dK��������ଽ������9�ף��6hZ���TI���m6`FM��5�k8�#�3��t��*$9d���oc�o��{m�N�;�/��(��$�����Ӹ�@�\��-�$L/'6l��tٚ�����3	ӑ�V�� �:��%J�][��W*)���?�Q�q5���.<���=Nݵ;ֺn]��O0qpw�X�ۋ1�.�z!\�d�,�u��=��Y�.3����B7wU΁�pH'D��%�_�0�ڴ � ����f!�f�����hdjӦ�e����XVK��Z�%ǌ�m�w��Kvq�Ӭ�n�߭<I�$���;uЬ8!Rw����>�����,̌�p���e�h���B7`b��f�p���y
6d�THYϓsm��ruݡxSf⣩�p�ܙ�����o��V��9�Ni7I���/_]�|�|�:���㇬r"w�ͮ�b73 &�c5�����`�D�{F�t2z�]�ۨ�N���pͣ,�W-u8n�U�J8j��CAc��13�pb�t�..0��M�!S�rн�jV��v��[�'<�V�2x��cͫ�$��|�좹A�@1��Q�P�Yn�$��ʲ�s�]r냦f��s�����o��^ul��gҿ(uwpA8��G3��w�^BX0f*���Br)�u�纲a�g=�D����wsB�9�
���'3x\J����@2������eg��"]�p�������<Ȱ�a��r���9^ݿllN0-�dݑ�髾MU�r�bs��$��F����6���bZ���jʉq#f֛�0b"�Q*���=L?	��0\9��o풹VQ!)sn��acr��Y���L΂F�8ҭ�����^׉�_�{�&)�Hu�
l�Q�_I����}6�y��T��+�E�]'�d9��9�c��L̅{Pe�FL�t0`�Ǻ/�}��	̜�����h*��3��\�Ϯ[�[���j&���3h)�9|t�z��ŵh�5ƿ'_��,�E%&z�"N�@mJ*H�<a�d�X�}���_��^�sb�2�iS��*/��ą�L�աa>I�������1H_0W�2�9�B�ni��K~�mZL���و�eb�@ڂ�͹z�%��p/q5�$7f.��߁��Z�(5I�-���U[�#�e�n����^M�ҋ9��,l�ȩp��e�뼮Id_��k�6�B��O��̺���}^�9.���"�~���-���a�Mx\��>��od�̫��'#M��/�S�q�����r�6��L�#՝D���X9n��E�3�}��fI�-��1��M���[W��|�I�G�[��XZn�un���ظ�T���g�.#1I�>��H,78�����r��O��}9/[5f�Ũ�X��˹�m�W6L�Ō�h���&��±��w�$��n>7���pb_]h���޺:�	N�ԭ����0Չy�%b�0r.$�Ss�qsNmN�[4��P�d�9 獷�*�~��j��O����f#'LB[����v�Є�c= ���d�EeyN�����3�S�f�_J�QX��*-��ڨ��L|Yt��1son��+Q�	��@	B�'L��,K�0\�����51��� զM��Y��W��X�	N��
9Z��w�6�Հ㺦\}���<��.�`؄J���ͦ6���$�^"����3�?3M}2k�L��׭���לM��E#���o�����s��23�.'j]�΍�f�vYtDNO.0����ùx�约H|�ʜIp��͸	��9`.��\w9�fVF�Cl��H�?)�:�s?L.�Ω��-��1x)��{�a8aJ\����:�
.�]�n�Tw���7 �M¿(uQ�;F/9"��$4ʖ�l�Ao���.L8�փ������3Wl�Y׳Jκ��&&��N+�N25���1�wy���O����n
���R�G1�M��od�O�'����a���|�RGf��i��Y>+	'�_����Zj�`�1S��e�:2fV���y�͚9-аI�y]7���e��p
g�f6� $Yy��t0�ΫY9�f��njbR�9��,��g&�ȹK��L��!&�<�E9����u9��.$��,C&s��́=<e��X+h!R��D��0�u�KyP}7� i�8!�(A� ��I�ë�>�pf�>��iU� Dm�� ���v�V� fj������ܺ>~E��q4෮In��(7ߺ�	S�
��z��d�?x-ա�u`���g�Մ)���]'s^����Ep��ོ�ii�9��<_�W����('<|�������D5�̍=P,?8@�n��Λ�\��_N`Ь�ꎭj��ߡz=�JT���*bB�*f�7�i9���A��5��nE��n��X��CO���[hV�:�$�Cs�n��-�:5j÷����hn��f�MA�K���lRNL��p��pX�/�5z�Sz�%��RGf�mv��c&��E��ì��`Ν�fA��	��dp$��w�zU���c�N�e�ޫ�v���5�8�/�!<��R�5d�����		ʢ3�λs�Bs�Ȅ���ZBg�j�y��0rnc�B��3FF�����������_x�D.�M�9�V��3x9ldY-ٕf��7G��\����{��,��0���V���H�0+p�؜ol�$������E�8��Ih~xQ#FM�'�E_��Df�2V&���X4cs�T��,��ؐ��z�͜�+`w�'��\�'�0ˡAw2=�2�VN���rsڮhE�)��,l'��$�6�F�����	\Er?R]��r���]эm���	�kG$4W�#'\elΪ{�漣�a{��iBc0�wg����,�÷�ųy7ɺs|ͬ�-
��9����٤,�UoY҇�%��E�Vs!�����s���ZO3pN��Cf٬3K�L�_ĺW�W��N��N��d�q��L�&��Z��qIb��\����,&bY��:4?�8h�u�x2�Qs�̐)�/�r���Ȩ��[��pf�QSd7�����Y#61�^�e�Q7k���m�^���8:���jN���j�7�J�L���R���fm�^kp��s���dݒ~V058\�"�r�s/b�=/]c9`�D�K9eF͊�YC�0�Gs±y�8n��Kg�Ѐ��&�Tf��z�S�X���0����uY��Of1�J����#�T�q��3��nS��,�@Y��w��	h*d����}���:�K��Ӽ��[���v?��Y�%3 �e�s��G �sr��F���
H�y�6��������X䠉^��"Pہ�
�/O�dY�˳0wa�9����>�jӦVs���mŜ��L��6�|���2�ҥ�Z�U��f�x 5#'��^����m,I�5�ĥ�3&�	W�zN�R~��|1�46�f�$�[�'�7`*�m�B���@�
�e��ꚙ��h���Y�ꠟ�;h�Yf��NN[�};Ho��Z�܄'�����_p��o��nc�lM�v���v��K�1P�朼b�lN2��;���PѨi�:�ͅ��Ixڤ5k��ըaC��|��˛�+1r?�4�6�R>/p�c&L�"�%f�<�����r3�z�%��e�9��Tˎ��z�-�ܣ	��c97]Ɔ�b?Њ�'��ͬ!7C�"��y���&���,�t`�e[�Yp���4�Nl&�R�^L�`�"-ρ��쫻�'�u��ەsPX����\�ȉX��3����Z�n̄)��uq��/9A�c�rc��Q�V2�N��Q����bҺ�!1�� �6{�P�n������x�,���)�_��;�N�#�XSz5jrhܰqfs]��+X��1е0`��(9��Ժ�&�5Iҝp�=En�T���p�$���]:a����)"g-��qBj;P�PA��	�, u1}��r?�Y7��nY�im��~�1h�,kY��Y����㫩��9ѷ$3hM�7�͈�����	�����h��ҋ�m�ս���j��5C���R9�'	�F���!ܘ�_�h�`�n��$���pg�����XW�Ss�GwC��0%_��,y7�7g�d��İhUݜ09�V4E7Z�*����a�T�'�ǹw$�/�f�6��L�\s��{�u�ZW��kg12�#'<��6��ϩQ�J�As��Iq������31@���tyo�,I������vC�nY�q���Ћ#I�(u�a8j�5GN��6�fn��Tj�9�ʺ��&&=2�h���f��n�psb<߉�L�T��R8}�ȉX��o�n�&Ѭ<�0�_���������mM_��Q���uZ��+	'�_��0O���ցJ�ꆋ��x�B}"g|�:1O�D���%�&���.� :r�ɜcs�U�f��a�!qԘ9l�[ͱ3�1�U�\�1*g�m/�Lx��f�����|/��T6+����QY��o�ܻ��&s�́�a�O�u��½�cINE����_��Q���p@�"N�@mJ*H�<a���:���sgy,�C�҆� X{��`�5K�����nNV��[��^p����l�8���V�B3h��[�K��Z��U_]1�8�#�f�3�M���f��`V�w$ZY�k<��kGMĪ�����7�F5]��^, �Ȍ7I�૶�g�2������mܰI֭ΐoy-71�X3��2����`\�z@�MM�B�)�a6jV��j���{d��6r����uOF�T��avi�Y�pEPsG��z��fbT<��T3�͔ݟU>�G,11|��AF���&b]��Bu5����dĄ'=�z��յ�Ӯ�ĊQ��v�Ir�9E�d�͸��-�d�σ�Ia�=���Y:]�P��|[g��Q����2sGՌd�ٲe�n��ښS�T�s	���r���ם�/DCfoSIj�y����aL�wP����Z���b��VS�_�df!1����[h|��3G�Ǧ�i��L>7���Y���-��j6s�s�MX�F(l�,��<���Pv������L=9�,���1uk}���q�O&F��Vs�9�:�op��#���A��Q83Қ8>ˋ̊8!�(A� ��I�U�4__.+r�_E0'�%g#��,�U#����s���ZL`6\��ą3Z��S���D4nN��<ǃ��c%ɠQ���9�4l�T���C�Y�j�,ǽ�\��2Sx���u�u��̙�f;9r�T�lf]6����ٿ�s3d�'։_��b��<�DJ�׭7��ƍW��²^v�3	�F�;��	 f5I��Խ`�<�Ժv�V�92�T�?�,�+}�3�Hᐹ���J����=!��Y)5jԄ%��,��u�{u��;���M�0͠YY5͵ըjn����M�9�8������~��YH�O��t� <�aA�9��bd䜨��b.�&ؠAsҞN̖��h���i�e���dn���2�X�j� 8>`��V�9�$O��[X��	Kj8K!]bBS�ܬ����$9�v>�Ac��[䇰-o���:7�5��fH�p9J����s�q���?ٌ3]���]�XB��ڰ9h7d�Y�C��9�&TR���eS�z�n���<��=)0��w�7}���?s7&�9�����#��Ws��_�`��p�V�$����qBj;P�PA��	�, k�<� s�s^�ڑvA�DO��Y���/��elf��r�W��O���ap��,7dF���:\�]M0�+<�.�E��m��y�44g��u�pbߐ�����9�F�D�g�k�%�����f`X�_�T�-�5^7`j�f��9y�$ү����4^�
��y���+Lug������M��H���~<5�$��h�sO��7u6����H��u���R,�uS�&b]�a���!�`���0�����S�Mu�"��p'D8�bQ�K��MU���~�o��aX>���[L��*b��'�nsp�	7lUq^�KvJ����i�>s�4���0�r���1u�e��7����R[�^#�Ɩ�ʬ���D+�[�E�{�<XXR�Vr��x���.�X/=d�����^n��,�W���9Dߊ�$�"�]�뾱!]��(uh�1�&�IV�Fcf����6���̀E��f��{bڲ�\�C��j��$�����M�!��w����~�o�M��İY�k�����]6d��C`4��f��0�i׷X�uY�F1p��3K���4j��)��v�����&Y@���.�B�y�����h+9�g��,�CȂv�Z����?��05z�ɵ'�F��^f&����}�#�)0��w`�����\��н�֖�n�����$�=�c��9蓑B��"�r��~�{lĄ��z/ϣ���H+��{� o'1ik� \��x�O�V��@6�+��-Jݺ�ѩ;����M�1���P^0�}�^@k������uX�l���[�M�죚�B��aC�рf�Wi�������@�x���jUV�\X35	����xΔ�[���Y5gK�_w4/���B^�v�љx���n	��Y751�D)s�F��b�nb�9��{��͔��w�[�5U�,����Gs����l�b��v�j�RR�Y��f_M�u`2�m�̙���2s���ssl���%Y���/�sHR�&Q��r�@�6����l"�I�{�z����D�RW� ���� �t?�և����y�w�ԑq��RKNC�M�sZ�E�&u���9��lz��U��@�qN�^'��{�ީ���|��Y�[��D-���ٸ�#�R#N���_�h+jb8��lEfeV�ML"Չ9�ȨY�3=&=0r��;,5�V�.����c�_��P�8o�Z��<��Y�m�����8/���?L�aC��uY�Ѝ�I�?���'���c��83�uk�9p%��\(d������`Ä�;���:ʉZ�ӟK{ɀ$�)�Y�n�ͦ�����x�M��!Y|�Y�	3�.lfb���Z`���l�Q41�9K�d�)��r\72rÊ��㈛�Efd;XF�K��Ԗ�A��	K����A3s���n����^�Z��"Pہ�
�/O�dY�����jt��9���s��,��˶�f-j`1n���\��0�F\߂|�O� B5`�;�!�0�+\�'�����Zw���,�CN°C�:�8��t���ܐRN���1v�E�%�A����h&ᣙK���0��:�>5d�LJ�uX�Ej�݀�������<��������^0ۨI��p���=KM�ՙ�_���ڼ��(�M��Lcry��5Q�^���͡e=�+�&���箠�ΰ�ZJn�p�� ��b��D��r��?��I
`���<]���X��͜�l��$M�asp�!7d��φ�`�ɬ�B^xj�4g�҅Q7���S����˃��SU?jWd)-L��Ɨtmḁ�.�a����q��I*�9+�yAS��8�I6u1�&1�����p��$k�-�O'Z!�+�fe���D+\�È�M�L���n%�T}��6�r��@l`�^6 �Z{N���J��$
9{��׾��`�f͗�m�M��ŰA�^b��]7+��`����/��z��Y��TG�_�ű��8I_�����J.c4hԄ�P'D���	�, h�}#�e�v�c�.k1r��VrjϚ�9K�5fv��pd���&Ġ��G\e����N��/\�uw�F�2ޢB���lf�6�&Y'g��Ydp��n��E)f�.~�nU�9������T��G���ݝ�]+3��U���;Ά$	��a����i�	)�y�l�����{NӅ�U�ݏ�����A�1�:�u�b����G��`����=h^��� ���.Yx���u�3�ۅ��}2,�+��"A�R?Ԥ�r�l�fܤΜw�����
/��9Ȯ�b��)v^�����t�T6�+��Z�{L��})��3��M���r���PR^�ê�����)�7�s��1�j�o]٨���'�=��w`�I')���tj�-�T���l�e~�]��K4�7so7���u�;<N�i��c�ޭ�i�T{A]39l.7b
���ݯ�~;���V�����Rk�M8���>����
1�8\*��U��uX�g�Tɬ�fo� Y��p�e�S؁��9B֍��G'5g�̜+FOf.�uV����z��Ѩ)16*F��S��d�f9T�[�Z5d��[N�t�<4WFLQ}����O��>�:_�s���M��:Ֆ/31�dƟ���+/͜jf���r�Y&)/7r`9|55���j��B'j/�28'6�J�F���Cs�%�Cۜ�%�c.�[2\��K�d�vj�#ktx5ǼTN���.��^qD��J_�Ac�p=Wd�.�T����Y尉��@���U�Sc,���v�WML���j������
��k#'&ƺ��8�ҳ���s⺉�h��'b�K~�N�ei&����8?+�ܾ�ą�|�����ʅu�W�4dS@�Ҡ�Z�c'�0lLlZ��
�/O�dY�i��k�vg�1�B�rj�}Z2���{ᛙpn��|�\�W?�k���Q�d2V".�3aI�9Ѥ��g�j.|��0�1Ӆh��9��O�Ό��s�:��Pĺ�㩴<�\�E��$?�WuٝJr�^w�܇s��Y���ey��o/�p�c9�d���9l\VB������s^��:��
&���ӰDX�M�9�Ԁi�+��Y�ج�ڲ9۪p��3.�?)٣��%��ͨ��'�3��>�Q{���t3KM׭쳜z#rJ���f�/��qs�G-,~3W���DFL�b����G^bF̡H́-Y8}p��Y��tS��砹���I��Bs�V�Z��g�طzI�E���f4Y]7`�Th��.�u=-�ތ�?�t��9-U�S��'�N2{pbذ��_�]`�����ܕk�&N���Ag�"���pf��4ኰx1f��������fb |3����[Y#,0d�,��l�p����a��_�I^E�;�ܐ��p3�U��?؝������H�.jNz7ST�P���s�8B��z�	S�h�[|WQ����"�"N�@mJ*H�<a�MS�.�Q����xN՞%f�Z��梁L����l����hb6�Wѯƍ��s�N]3)K�a.M7hԀas����?ho�&�p��<�2X�`J��T��2^J)"_xA8�nU��)j��ir4����Y�l�s�_���E8g�uY�a������و�R�&���86I�?�y�nb�N���-Wnm���$*��m8g�:�)��Y�+r6m	&����f���1�^��8�����՗�jUn�I9��&F���`���ب������@ޠ���pޱ������
>�//9����p�:��լ}���s�n�R���pd�ֻqc��g�T΢F�&	 ��֨��l֦Rv!�_G��jb9d���T��̻�\�3��$j�u�Ԣ&�1�%����~*��7I"��-+��o��ꫛ~�.,�$@D*\�IcӵL:��
�H��I�X�Er¯̀�ԭB���mI�ϋ]'6n�D��@Bf���m�p<r�͑ٔ�a63Kjf4�/�f.��53n*��ʺ��":��$��ꊹSf��rsU��9�OL5q�/�r�j����}=���|�f-S2d̈I%uO��Y�3Q�ʛX�g��(C�י9�B������8!�P�p1�`5��AcϢԝ��3��������\�݀a�� F�Q�P�ӹxT��Q�0���{!��MXbDeÚ�Y���L-T�	��@	B�'L��������x���C̒Y���{�<��_���4k1��pY6f�@9���
�ob�Y'6����ج�ǹ$�+\�n���VLa�����,%2Mx1�n9/�Æ.�j���b^2딬3s����m	�DXNhF��j_|4�T���9�)�Kw�PH�ΠI�Xy7l���ֵ�+Θչ�a*T���1��G�6)�F-ؿ=K��%-�3�q~�[3���aFN��./4�py��5Q�^����t��+�&���ҒES��N��Rr'��=�7I�l.5��1���&��y
f�n���W��ɬS�&h�ǡ嬦��f𻌷�#GL�6��z�AsfCsk���+�py���c/����`��f�E#قtH�p'b]f��-�\�B&<�O���uF�F���
`�P��&
Ŭ�7��i��F8Z6�-�� ����/F͉�f��p$R�aэ�xS��$�9%����M>��8</���ab��+h���^{4b�D#goݖ��^-U2��Jf]�6F�b�ܠ˺`W��:�HS&�h�k��{�ذ��,�́!��#N�ףga���5a(T�	��@	B�'L����(�0\����r��Kjk��<��sX>͔�3��]�%�|�TV��ד̑�R}����f�[+n�L��n�z�[�5�pc�#敫V�k�l���/�T(�[�b&�ډaSa3�{��Iȹ��^Hќ��l
�V^̏��L�����p㷢eY�9��!4&��]���v��8ò���IƸƋs���Jµg3���Ȝ�	V/�M�7�M��.�-^�K+�����ݱ�&�Z8oQs���*�≷�hԌ�I�܀9]Ь��R�f��j�nb *
M�F�Ã.+���6K����"�sk&gmϩ�V�:5�{��.���氺L�,��#&D
��7, ���d�2}�ێFL��ШQ��U�F5Y/\���sJ�K�2�I.'��:�Y�� v�j��^35KG�6	?#չY��^��
M:�fa��h�S�n}��>.%7��G3�_��+JF�Z�Pvq۪�,��y4dj3�輊B�W�]Ĭ�m]��}=�T͏��%��H�'RႽ8Ѩ�c�̕I���w�ρ�����\�jVe3p�A`6\����R8��0���u[0ج�F�T�O�S~���1�(<-z9G��EV�<aԬ����4/d�,�p2�.ܿ*b�⊼'��eg�_�b)]x�_w5�])����r��@!��+,��a���p!ZhB3j�)����̗�¬�ޚ�Q�͹u-ጭ��&�1I��_�3Z��(�M���B��z����P��8�.�Em��W�Yb�t���M�bN�u]�[M�M-<H����2p�x=(�������]���so"��H�9nv�%��m����3���z.7r�$7J�Z��?��$��CZ��S�8�݁+�-������en�D-��nwq�\t9a�1������jԀ�lX�42nܸY��_dhؘ�S#���_-1g�FV�M�
���Y3���wQۿ;�Lxl���f�FM�΍���;���H�pg��D-�<\f��r:�̈́+Ff���p�|�ܕ"�"N�@mJ*H�<a����� �e$=��֕\"gR����4wW��6�e9/��gu�AS��&[�YvnN�T�uX,W���L�P
]7��ʋ)��I3r>G��lغ�1�3�/17��+�|����:3�?`�ݖp:µ�C�:�RD��H:ŷ30؅h^�ľ3)�ׁ����ֵp�e�e&A�������e~��$|�Vxڌ=K��%-p\�=5ck*��}7f䤨x��ջ����U�0�ux�=6٬��p�8v�����+�ġ[���&N pn�"9�ѐqST_s2�Gr�@�����)/�A?�k&I4ͺ;�jj��h��f������ͩ�^d�\��/�:���+�p!۬��@��v�/lKi�����P|I�v�p"�e6��9q����?�����), h���D���t��|8���nZ�pn�~�8�
ᬼ�e��!RH��>����@���WC��������l�CN�5���0J*x���n�<2�FL�(��G���/�Zy4�⹹61������]i�t��ʲ!���Y�uZ�b�fQ���O��рY!I_�����J.c4hԄ�P'D��%�_�0�r�����Ŝ�k���,����ڳ�`��5fNz fjh0��R6�:��YWld�$\{���8�Rxx[S4��j$Y}1c��<��)�É�311�; @��Y��bsޭԚ/����
O#5�7�3�Mҙh�ˎ����8g�BO�Ź�4n�,�c?�~`η� d�9�%2\�,��f`��6ဠu��J�_K���O�M�Y���YL������-\����ZhĀI���t_��uvs�^se����Y��9|��9��>x�9$j!��x�SM
1/\�n���J�	1^��k�\ɀ���pH^�N�CJ��:37h�K[�i|4��ـI�m�B7�M��>��D,dΘ���X�����q1nj�f���#{�q��oz������f�ܫ�,<��iu_����%+ᬏ8I�]X�_�}l��Z�1Af!��j2�S�[�j�\㩬θ9���L*�C���Q�F�2�ST(���lаI-�T8�_�Es=�,e7IЋTh�D:O=9I_7s��!我�i��]�����^�58N�S�
o�p��.8Iգ��#�M.�(<,��;ky?���cfX��;�$��,�C݋���he�sҐA�bVb�ZanĈ�Θ9yټ��O�*�9�O�C
����
��Q�f�l&&4ï[�\*��1#��Y:k M�^�㢯$��
��p��h� �&,1��e	-�:��9�]j7�d�4����w�I�E+���p8L�N���c�"��>�aG��h�Æ���&ja����u7�Bܠ	W��-����b
|�/G��?����p�Q��7�F51L�Rx��Bf�+��f�{'�7�l3+y����8�����w���Z�`�AqKq�MXbD��n�-W9>qBj;P�PA��	��M�R0�q*�9���Y����JN�YއR2�K���BofB��r�:��\q7d�~6\���Ñ��n�`"׽cIlv]�l�����忁e�zݡP���Yt������[�hι+�k����lT͹�b�Kp��sr��~n~��bS���D��U`s���ғ��f��D5pN6	?#���ͰYt�z'�ґ��^����4��L�q)�kJ�u_^��tAs���
y�Y�O�ͯ~������Y V��輊B3`B�.��0���t�8��0���KM��V�:?����.�u�<�[&Ɂ��q��g�2l*i6�F�e��'
����2�C���w�5��˓M�G6I��x�e=��%H�N����*1^��<��w��B`3�Y3F7p�U� ��T������
�L6h��2�Wg�3p5�ȩ�c��#湓X; �9��EL��" 0df۬���&\1n�0'�1ّ�q���Q7q�W��,Α����9���$7t�n�:�����6'�ڜ+w]X%��۲�^�;�xo��t�Oi3f֙LL!�琤f��-��R�13}+rfD����uz 5\i8�H���,��s|��S�7u�0#'Y�ܷ��AZ�e3����D�V��O��u3�I8�P��}��S�p�l6r�*�n~��,��_4/ ��`~�V�8c��_c4bb���� �d��B3�u�Ĭm��o�	�\���a�6rl8��b����2>S٘��Kh�9�Lk�^hV�a*ń�P'D��%�_�0�Z^����vKq�,#1'��X{�x�%�jd��]4@�Tז�1��C�5{h8WF��T�T'��S-�V�M�h��2e�l�u1!S8�� �Y�/ɺ�u�Y�hr]w�<�7��հIש}�]�E��L�pap�&4	����U`#f��(���r��,�f�$��Tw�-�C�8'9��5���{s��dp�[3�_=3j�ڋAS�|������O�8b*����G�U��0XM�.�-�C���Ա.�j�f�]��
�h�����ɩb��hG�Vl�6�l�2#f�S��lW�@�Q1�����:��Թ�x�^��vb�t=Wz��l_uPV6�z��IB����?��Ʉ�b�K��)���D_����T��@2�e��1��LJ6\Vnٝ�+�f5ݔKe���?�>/���ŭ]�R���2h�喌���y��l��Zx�-��Xc�R�[�%���\Q�pw�^��NS��bN��L���Z�qgE��I^7+��RN�y�	�rdbʖ�Au�-ǫR�~���󢹀��\������B�3ny����H��1�9�<�J��L�o�!�$��u)_��L-<�Ͱ9���֓�6��]�� �G�T�S�D�0Z+9�H�&Ɇ�����-��<�1��\�s\�*��ꦀ���a]����/0�1S%��l�s�[2pȤ�x�_�p��>�c�G�g��,#f��oo�L-<]��݈����9�r�T�@��/�Պ�E��p��[-����M���B�E���"�e��q~��|]�3�F�)Py�8?ù��5\���rY���f�4ܰ��)M^����]}4a!��y2/�ϊ�n�g�,gy�bR�q3t��̀)4Y�uY祳�r�ւy��C��.�]��l8<�I��d���T��l7��� 710�zd�4���?�2���Q��.Dn�o2g��������\�$��,2���K�h=@�1V�nEbJ��]ټV��ϺjV�D�ೖh�ke���V��f��S
�Z��rO2��UP��~��Q��8�7�t��Hwo��22�FNv�̵�N�r�N͡�鏝U*:-���o!\LM�F��}�4hj2��F��&���.h1�g�Zz4ɹ`n_����9����5g��Mc�>�ͺ�Q�&�8ϖ���1�@�$؜~��ȅ�������P�9}��U'��#&�5�Y�"w�����[�C_L87u�Z�6L���l�z	�Y ����R_åt��Ʌ��k�7����7�jl���2oC����-��H8s�φ\L�Q��A��@,7b&�S.f6-@	B�'L���i*� s�?�@�����1���ej�~�E����P���^�ln�29�]��0�n�w��������S��e3S���y	�f]S�ZW3j�=��;�����s#rV���U%16�~�M�Դ�b��Y��q���*����֬ˉ����0%�����!g@�e~����:']׃��\xըq��O����М�j����W�@���Y�g[����R� -�%���������5gT
��1{3�,i4Sv��i:�05|=P��H�\X�o�]f�\i2b�	�L��a�]?������b���s�̹���S[v����`d�$	y�����l�.��e������%`f�]7`�Tد�-���][3b
̬��_���i���G(���N�!�'�c�f����0�}�÷��_34q�[�h�[T�E�ˈY�`�l��M��/�Q���y�W��F��ܬ{dnf���s�:��G\~K�̹�&<e����H�#��edƃ� ���439�,���2��f�g쓉�w�՜nVSLU'B]�Αd,S5hЄ'}���%�7s�g�U�	��@	B�'L�6�4���嵚W�ɴ��r�YB`��N/= f&�
�#�A�R�Y���pnfu7�lѐ�6G+[�뷙#�A-o7��5����#�f]Ѡz�Ib~ѡ��F͡bu��~n�C�pA%�9����]`+нbM��±"r���京�&� �f���U��ɛ�-Jي�N��ݾw	�7����A��B��J8r���$���R#C�=u右��)&�mT�f%�w����(�[�c��&�]�c\e��É��uWs�.��[ǰ�-/7G���|֪Y��4g�!�z��ӏ��MN3wN�4Qff�'��l	�&�sd�d�lR>�N�e ���ঐ������h�W��!N���V�@�{} �nq?�1�m�$��R���w|ހ�uw�z�ۦn��m�����?�K���W���u���3Ӵ^�`�)�&��7���bN���s'<8�bQ�;��MUo��|��M�whZ�5 ��1�Vqskp��!I�u?L�n���ѾxCd��I��������X`�n{9��Sg�R�|ɜ rZ�8�O�"�}��sI�n�p��eN�Ϣ�=>,,�O���uD����� G��ub�ˍ���C����8�b�M�
�,K7j�m�d	�#ա9��cUL��y�PYN�p��wY�zi�����i��\@�ά1I-�{�ᵭ|~�%r
/�M��ւ��Y7��7�Ь�
>�-�`�J���N����9��!����bI�x��<�5��qBj;P�PA��	�, �hy��˲s�,��.FΒ�3�L��Y�C���l0S���fG��atY��r��vn�T�R���f��4I��7hZG$3.r؜�f�ل�/�E��#�a��7��T�5�d���7p�u�x9��+L�fl�r�&���^���5�l�Op6vdRC�li���:t���<>�����&�-��1S1�1���?)�ՙ9�1G��o��?��\0��7u)n �biSs�Vӷ�&[�W4C�K�����u�K�л<����������7t�l��{j�rؤ�z�2yB7�u�t݂��dN��KN��b����lP?��f��]���Ш�+h��q��4[�}��1b
�k�Z9-wjx��s�$#�'�Sk��]2n��i��݁$1W�6�m��Yؗ��*�u!�����pȄ)92��p�+F�J�C��q�fт���ew|�1cFN��������^������Yգz��I��l��3h�'!Q���98���S���}21�.7bĨ9��Tu"�e�N37RjȠ	G�h�!�x6��?ˋ̊8!�#I�0m��@�
�,(A� ��I�����v+f��͂���
YM5�s�-@�g�r��@���M�2�~76t���.���lF�PLM&��r�%<��prY�nq�9����X��!;�sw����)�榭�K�\�Wl'K�J̀�0+�f��r�s��pмK�nM՜'h
�c�Bu֫9^ԈQ�LTU"ԉ�un�C�]���E^�'����D����W�f�w%ύÛ�D���Ds����pU�9,�kgfm�c�ʢ� �a��f���B���f&�R�^�rĘs�k�*��R_���d��2�q�q�Y����v�=��uX�
�s�^�fP*�˫�� q�c���1�fy|��V��.��{�$�/�s æ�=&�����8]ΛսK+d꾫و�e����I��Y9�g٪Y�`*S�\�ź�Q� ��q$�Q3��&�n�֗�9`FD5�)Z��X̀c� qۦfQ.����-�g[8����>��YI3l�߮cÅ�2?������Cs�7��6~�����2��j�I2!Rf�O��vM݄ɿ��0��
1�L�WS��ۇ�
!Qd�х�f`}5�ܥШ	��ֽ�d�
R!��7�C��f&.�Y�kk���MC���������u_�eu�A��i�|[�q*��M��uG3�n����yY��}h�Ӛ�:5`��I���u�?6V9��mh؄'�B�.b������l~srn���Z�$#�J���O�ni���揙��lܬ@0�r�l��[�3��>�K�&i<�%�ͽ^ ň�XW�C3��44���'����9��t��51�991u�Z��ޕ_�l����X�)���$><��ډi�-�{r���&�?|��Q�l�:8`�ȁu�c�6л�_kq�&�eŖ������%T��� �&b]��U:����D�+�Ł�mrƐv��1��N��N�����9��
^?U���R�~8fF���ߺ���B7���H�O��zV��A��}�,U/Z��]·:6�C�R��ԉ9K��vnơD�3_�aAΐ\��9���Y�QON�O2dZ��v�˙��#gt?�Og9)B���3�i��r�A3�X��=������fc`Ԭx�Y��uy/�;	'�R�5b��oj�y��g�i���<|��^�r7�kԕ��B_���O�{���E ��ЕW�^�y��ON�['D��%�_�0�r�������@�B\92KdAV�=��
bv7��Ќf&��id�Q0gթ���k|XF�M6���&���\����:7b4���ܜ��pM�B2)�����]��/J��⦟}pRGsِ��Y=4fr]4�#Ե�~���[pԄ)=��!oCˬ��93/^�fR�G+�jx����Gs=��b�j7P�W�F�iT�;8C�&Eg�:4�ޡW�Ɂ&!42.n���)csX[�O:�e�X�c�����;F�R/���o�}����V�������%Y}0X�j�dV}���2�� �WΥ�a��[��Z��2�7��n���Ò�b�Y�pNҕt�ם�������m��Κ�ܙt��]33u}Р�S��]�'GL��g��f�E��fɬ۹�4�$��R����r��v�KA:��`6���:d��9I'��X�u_e1d�l�P�	��A�S��4S�����y~��KC�uYDk�F�T��-���Sϼ����z1��Qn&ze!����ᐑ�&<�է�j�9`���&<����@����T��Рq3�����(���f-WbŲ�qBj;P�PA��	�, d�~��W�������A@���y�aα|�n��	,����<��qg	,�5[�M,�54����DC7gh��@��Y�Ճ�&<u��Ԇ�w�Mĺ���Y�N�:�i�����.�-�S���<�9��̤E(�����f�l��%X���ꉉ�C�J1Y�ey���-74���|¯���1F���ck�W(�C�3j�$Hq��-��b5�Nx*�q8�%;Q�D.,^���F��3�����f��IP��{}�����u[R	_��-r���?ЫI��PI�Xa3�5-G�pkKԱ��b&������c�h.����5X�us�{����V{�텇g�a1/�Si�.31j�R-uFb �ƥ�2�V�f����.��ݒ���$��Rw�~��Xޥl1mlQ�/dÆMh�E�+�lBˈ��"�Ko�yc8x�.���e����(��"�g��C�2?�-ة�n@6h��Ɨ5U��B�|X4Ko������Yv�/J]8�f��&fwk�FL�T��81�F�尵����FW�r)��Q��a��E�挃s���a�J37���Y?4S��̀Y9#�Z���l��lzE�㦵?�nJ���^�6�:1�N͉Hf��/�F�
X����O����'4�$�����h��ZKa	�Ca�W���B����M�Y�%
&,<[w9`)�u\����v���g�I�h3r��}[7]�)3�
4)���L\B�ON���c	6�:4lN�ņ�\"��H��p��L�����lO���<Q���m3\Ȱ��\��݅2��r��\�'Q	g�|�'D*��E��[��*nR!��z����lE#&D�X5+ε4�&<��@�·5���1@�TW6=�l�&D��L�ORy]��᪬8v9�����"Y��"+��N1d�99+g���[�1s�`3�]\�R���NN9RH��j,������L�*�,�Ņf��0�.�*�V��3rԨ9�ޭ��K`�Wga:��LKX*�8I.�8��)~G����y0;֝c������/x���5�v7�M�n���Y����D��J�1��^�23!R�[1��5����*����f!��hݸI�y��Ž�͒���S��dؘYg2�1��U�y��፣A���/��-?�3t�R}�fcl�̏Xy]�,�ͳAcf�b��T���1�11�ڽK�+0=9��ʕ�*}pAZ�q�
6�h�,\n�:��.P��� �Q���}-C�2��Q�{e��f��<�@71�10�.<���f�d�5a33l̬�	�}%��-3k.�����I��Nn�ٕ>)�T����Z�II0�j�ϝ�%j*4�y��~��q܄�r��N���� �2�p��rY�cc�ɘ	��pj��Zf�\R9�)#����T�p�N1{f�Ւc�=L�UsӅp�wsg4jĤ�܅g���q@�J9hȸy�5]�b��H�r1�k0�s(��ʰ�N���uYQ7�v��aA]�����\��F��pd����B�'4��A����a�8v�&lԌPͼ��F�7rB�2L�~��094�R�����3+�tZ�w���As(p� �W��sJ��1�hƅ��k���M�n�~Y�Ÿq2S�&��8Y�k�&Q��+�8�щ�d�li��s����,卺i.R8j�v�u��l|�͘Iԭ�1a̏+�u�)r��l�L��Xtp��J19������&�ߕ����Qqܿ�+�f�,�T���6zܩA�^��k��$�R3<����q�e0I��ܯ�tgU�g���-����lz3��S}����rVhW.[8Wf�V��
2�+���Ҝߓ憊�2�r��eI�v��)V�^�Enf�/�U8ߦr%Ќ"`�\�\fǂ�Rr�k���Vb3jF�xf���MSrY�'��y8nJ�Sr=�!���:���0*f���vɺ;�0��}���N{0��ˉsb	,��/fҫ	�^Q*�K9������u]ńLetF��Č�����&YkNfZ~��yw/�l�l8pV���s�m�٬�V��L5�F�(1l6�Mv =R�Ⱥ���vL��E�g�K�;�$*Ō�d���#&l�g��t��d"W��'�3��Е���'X�1L�R�f�oj6������rْAC�-��Q�����T���o�J1��g�����F͠xY��P��͑�p*�.<@rp_�p�骳	F�iA6��&ܬ���um5���eZJ�6`Z�͸s�_,��/'<����=4��$��r��Ƶ#�i47$�:�Y��~4UO9f����2f�~���P������+��G3�$�7��Z�����لGPk~�fͬ��0�E���͒9H_���|��8!db���-�jԬ 9+`cB3c��YVwi��=57bѓq���	[�Wr!�S\�}1���C	({�x9ۺ9�r�?��{3G[��/���}���}=�����9�%!�Vod�.��#�1N�Gf��NO21����\�-��

c庮�b��Q5a�y��^�}0a�|�b����Q}1)^$1f.7�9����~>,�U!�$��Mx�}��ށ������r����e����kF�+�ң3<eiA8jVf�L�s-�M�Y�K�LRț�s�^�k�:6��E�ʹ)�Y�sA�"��F��Հ"��s�,;3�����	S�Bp&.V2��M�����C����9Qg澉�K��u�>��1���O���T:�����KĠ��u��yh�"0dԌ�`�I��ns|�	W�?�Ϫ�؄ɟ54cf��20p�dI#�۠�hjT�X!\���k���y�).�Y~�6{����Yy1#�e �b��5_�wH��IԹY�%���w@0<u��g���,�KnVS�'�X������r�O�[�8���7i�*���pd�j�T��nl8�y%�D�-
|�Ar��F�����v��i�asW���MR�u���}�W]3rB�nYk��5��(ur�,�pܰY��&'A��n�]�5����@�vh��I֩�d�^�l�����N[1][4f��'�9��e���PNq�̄X\k 'Luэ�RU~0�5Z����
�!P�����b�H�S�Vo�Mw�qfA{���c�&Y���'Y6h�l����q�I_w9�fe/��E �B
�Mn~�ס���������o��Clb���Hu�dwu��|�ܠ	O�!̀�\�0��5�����_�j#�4[�j��ͮ����ТA��ͻٌ��,��"N�@�����&Y@���>*`_4K�>��rJϢZ������3�/l�y6֊޻*�R�Nkx�٤p�nɞ�~[@��ԝ~��uڌ����2l^�9p�l0T��gF�����&������^��J!ŧ��e������8cS!|ۅy��^L��ԭ�	w$<���ubj����� ���´��A�M��̌����
�M¿(u��@8�]Q3f飸��#�*�Q�&Y��ت⏜w��[[5�HzXm1g�ڭ\W�ׂ���ٗ'<u��TY�.��OL.Ss��&�\Tl�o׺��F��_Q���xyI�_���ΆͲ�����0_���f���$�^D�jlt}��[N@f�N��F�3��L�#d�fV,��͂�f%������JkzF�l��(�FЬ�JȉX��u����lC��ύU3��,32ap�ub��s�j��`5�Iɰ9�A���:6`�\H�w4�)򯂘���2��{��_�ur�@�������S]M&Q��h,�V��r ���ltшIZ�1�~�Y�;c�}ɝIk�:�fFg˻�:-90KL�_{3`�d�Ɍ�ItN04h��ǩC�,��i1�v?k#Ձ��E�<�^8��0�_8мbSk��L�ܿݫ��a�b�`|�[1+�>bܘS�?̯�ڭ��� �◝s���)��v�����&Y��3@���-��k�8p.O�9����n�^
�c�r*MN3�x��&��ח��3sj�	Sݪx��n��Q���Α'%��w����]�.;��1Ԡ�Rm�,�nĨ�s�2n_"f�h���<�P�9�V�N�����I3oH��z�����Q��廘Vf2`؄ɯ��n��لɢgS�2�c�GRGL�m��uaY�V���7K���%����y�a�͢h2��J�As�jr.�%x�^F�d&<u+��:��W5r���A{��C66a�[�������B�f��n�v��*���]\�TM��V��*������E��S;���s��A��y���y���9	yЬ�A�0�h����_C1h2c�������Q30�u��Z�Y�d��������\��$4�V�>����~���`�8nJ�hq�\��o+�f�[��C��u����։Iɺ�M�KiɆ�*Q�Ӄ�q�p˚����mr�q�|��uYhKmi���+L��V��21������67��_���w���I�wp g�N�o�mbAs��+�D����F�9��T�@�\�3AN��Q�N�b��#4	����Y��4o~Y&	������,*2p*�¹�jj��X㯙��R#�9���Z��]�b,����It4t��a�uD'�^jb޶��N&"�J�RY>7�{��� �K?Ā�����2�#���a�i���Yw7�0��Dh�-��<.��'Yw��̀�1fB�.�fN��v��@N"ׅC�x�B�np��u&�D�Q-�eA�*��M>�5b�D���u�Ee�e�=��!9�"ul6��9T�*��)�em�̲W�U�ԭ��=2�ﺦu��`.g�5KN��m�@�<�$���
ug��:��n�g�b�;�䨑ua��Z��x�ȸQ�0�y���5�è��WsN�.�Y�.�_f�T��cSp�ےI֙Y��o���qS�����pbj�����������3�����,{�
���mѰ�XW|C�<o�J-8aJ������_��8`V��f��,'Lu�$g���l������V'���dz5f���hV�Z�)de3���0Ia]%3'�1n�r׉��k��Ԅ���R|b3+)NM]o	���cR�S��mUf��y��nܸ� �D�a�Qt��&W����IE���i�`��E�[(��sa�_���Ә��u߯�Bz6Hd��aeo�:���g�٫f��9�'��C�5�ۛ��P,���&Y��lƯU�C]w��9����H�����SM׹V��-ϋ&Yw��;�V��y���u9��6[�I�,3냦��*�9X�9�&�V��M��Bt�E�K��2Ǒ0�_���J5��8;R7K�0�ɹ�����E�;�7w0]���H�p����8�eS9��Y���$2I����C3�]`j�Z�-D��D���r��~dj�-�g1给D������]��/ѻ��I��n� 1fI��߂���AQNR�(ur�p���,�uv��w|.�3��J�I�тt�y��@��Č|+�J�IB�&Wj�c�T�hu�?5��w�{�%����8Cp5�N�bX��h�l)��v�����&Y@��>�,L`���Pl�lu���)=�b�؀9AV�L+f���>�
c�a�5���܌�;�^|ǝ�!ש�.G
���QuQ��b��P3h9�} �s��&ݥ%��j�v2+�Lxl>p� 3dkl�d�r��wL�C�Z��&��d��q�։�
�r��I�̻ɴ{�f⇁Ӿ-C19�i
��vd��M;��T��fٲ9��P��{��ʲ�2a��G�ALc��,"6wN�z_��_��XP���5�k�����KA�u+T̑�mMQ�H6�T���:f࠹_��A&L|30�"�c=Ȅ����܍C��
ćb�GsީYp���kӢn���Ϳ�Mvi�齃�H��L�������b��:?��guu���.���˩|��(jΦ�O�{��2+�����j��K��� Sw�~��Ǩ����B��6su���K�̪<T��������I�M��3� �9nn�e�����9U�DSOLJ�����artOz9���us���@��f�9x�ӊ�	��}������bƺp�w`#s�l�~jԄ���-c��W#f�l2n��� /O7I�����rt	S�ʒC�'z��F�#Rsm�h��--===== CDL4 =====BM       6  (   `   `                     �       �    �  ��    � � �  �� ��� ��� �    �   �    � � �  �� ��� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� �@� �@� �@� �@� @@�  @� � � � � � � � � @ �   � ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� �@� �@� �@� �@� @@�  @� � � � � � � � � @ �   � ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� �@� �@� �@� �@� @@�  @� � � � � � � � � @ �   � ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� ��� ��� ��� ��� @��  �� �@� �@� �@� �@� @@�  @� � � � � � � � � @ �   � ��@ ��@ ��@ ��@ @�@  �@ ��@ ��@ ��@ ��@ @�@  �@ ��@ ��@ ��@ ��@ @�@  �@ ��@ ��@ ��@ ��@ @�@  �@ �@@ �@@ �@@ �@@ @@@  @@ � @ � @ � @ � @ @ @   @ ��  ��  ��  ��  @�   �  ��  ��  ��  ��  @�   �  ��  ��  ��  ��  @�   �  ��  ��  ��  ��  @�   �  �@  �@  �@  �@  @@   @  �   �   �   �   @                                                                                                                                        gggggggggggg               rrrrrrrrrrrr            '''''''''''         hhhhhhhhhhhh""""""""""""hhhhhhhhhhhh""""""""""""                                 ������������||||||||||||											||||||||||||������������												   																								      hhhhhhhhhhhh             JJJJJJJJJJJJtttttttttttt     ����������������������     ,,,,,,,,,,,,||||||||||||           tttttttttttt||||||||||||tttttttttttttttttttttttt                           												hhhhhhhhhhh            												tttttttttttttttttttttttt                                                  ������������������ ��������� ���� �����  ����     ������� �� ��� �������������������� �� ��������  ��  �� ��������� �� ��� �� ���� ����������������� ������� �� �� �� �������������   ���������������������������������            �����������            JJJJJJJJJJJ           JJJJJJJJJJJ           hhhhhhhhhhh           JJJJJJJJJJJ                            hhhhhhhhhhh           hhhhhhhhhhh           hhhhhhhhhhh           hhhhhhhhhhh                      hhhhhhhhhhh                hhhhhhhhhhh   hhhhhhhhhhh       |||||||||||             hhhhhhhhhhh											�����������           											hhhhhhhhhhh											�����������           																						           											hhhhhhhhhhh											                      											              											hhhhhhhhhhh											hhhhhhhhhhhhhhhhhhhhhh           											hhhhhhhhhhh											JJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJJ   hhhhhhhhhhh											 mmmmmmmmmmmhhhhhhhhhhh											|||||||||||hhhhhhhhhhh																						hhhhhhhhhhh											 hhhhhhhhhhh											'''''''''''hhhhhhhhhhh											'''''''''''hhhhhhhhhhh											                                                               ����   ���� ����  ���  �����   ���� ���� ������������������������� ��� ��� ��   ��� �� ����  ����� ����������������� ��  ����������� ���� ���� ����  �����������----------GDLN 10
6438 0.0000000 0 1
7000 1.5707963 0 1
7586 1.5707963 0 1
3358 0.0000000 0 1
751 0.0000000 0 1
9091 1.5707963 0 1
10783 1.5707963 0 1
9771 0.0000000 0 1
478 1.5707963 0 1
1001 1.5707963 0 1
             CDL3����\C ����PVBM����6(  ����GDLN0����   ������������h$1��1$h